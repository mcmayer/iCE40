-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2016.02.27810

-- Build Date:         Jan 28 2016 18:04:01

-- File Generated:     Jun 5 2016 21:32:20

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "uart_top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of uart_top
entity uart_top is
port (
    LED_o : out std_logic_vector(7 downto 0);
    RS232_TX_o : in std_logic;
    CLK_i : in std_logic;
    RSTn_i : in std_logic;
    RS232_RX_i : in std_logic);
end uart_top;

-- Architecture of uart_top
-- View name is \INTERFACE\
architecture \INTERFACE\ of uart_top is

signal \N__3943\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3931\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3922\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3859\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3841\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3829\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3779\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3747\ : std_logic;
signal \N__3744\ : std_logic;
signal \N__3741\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3717\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3715\ : std_logic;
signal \N__3714\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3660\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3654\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3646\ : std_logic;
signal \N__3645\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3618\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3612\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3577\ : std_logic;
signal \N__3574\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3567\ : std_logic;
signal \N__3564\ : std_logic;
signal \N__3561\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3558\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3555\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3537\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3531\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3527\ : std_logic;
signal \N__3522\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3513\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3501\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3451\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3447\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3441\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3439\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3436\ : std_logic;
signal \N__3429\ : std_logic;
signal \N__3424\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3419\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3391\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3363\ : std_logic;
signal \N__3362\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3360\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3354\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3310\ : std_logic;
signal \N__3307\ : std_logic;
signal \N__3306\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3304\ : std_logic;
signal \N__3303\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3301\ : std_logic;
signal \N__3300\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3298\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3287\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3282\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3274\ : std_logic;
signal \N__3273\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3271\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3209\ : std_logic;
signal \N__3190\ : std_logic;
signal \N__3189\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3185\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3178\ : std_logic;
signal \N__3175\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3169\ : std_logic;
signal \N__3166\ : std_logic;
signal \N__3163\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3157\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3123\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3104\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3090\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3083\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3067\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3036\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3024\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3013\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__3001\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2977\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2970\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2967\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2964\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2932\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2920\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2911\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2898\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2896\ : std_logic;
signal \N__2895\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2890\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2887\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2868\ : std_logic;
signal \N__2865\ : std_logic;
signal \N__2864\ : std_logic;
signal \N__2863\ : std_logic;
signal \N__2862\ : std_logic;
signal \N__2859\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2851\ : std_logic;
signal \N__2848\ : std_logic;
signal \N__2845\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2839\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2823\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2788\ : std_logic;
signal \N__2785\ : std_logic;
signal \N__2782\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2779\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2772\ : std_logic;
signal \N__2769\ : std_logic;
signal \N__2768\ : std_logic;
signal \N__2763\ : std_logic;
signal \N__2760\ : std_logic;
signal \N__2757\ : std_logic;
signal \N__2754\ : std_logic;
signal \N__2751\ : std_logic;
signal \N__2748\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2736\ : std_logic;
signal \N__2725\ : std_logic;
signal \N__2722\ : std_logic;
signal \N__2719\ : std_logic;
signal \N__2716\ : std_logic;
signal \N__2713\ : std_logic;
signal \N__2710\ : std_logic;
signal \N__2707\ : std_logic;
signal \N__2704\ : std_logic;
signal \N__2701\ : std_logic;
signal \N__2700\ : std_logic;
signal \N__2699\ : std_logic;
signal \N__2698\ : std_logic;
signal \N__2697\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2690\ : std_logic;
signal \N__2689\ : std_logic;
signal \N__2688\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2686\ : std_logic;
signal \N__2685\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2678\ : std_logic;
signal \N__2677\ : std_logic;
signal \N__2676\ : std_logic;
signal \N__2673\ : std_logic;
signal \N__2662\ : std_logic;
signal \N__2653\ : std_logic;
signal \N__2650\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2642\ : std_logic;
signal \N__2637\ : std_logic;
signal \N__2634\ : std_logic;
signal \N__2633\ : std_logic;
signal \N__2632\ : std_logic;
signal \N__2627\ : std_logic;
signal \N__2624\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2613\ : std_logic;
signal \N__2608\ : std_logic;
signal \N__2599\ : std_logic;
signal \N__2596\ : std_logic;
signal \N__2593\ : std_logic;
signal \N__2592\ : std_logic;
signal \N__2589\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2585\ : std_logic;
signal \N__2582\ : std_logic;
signal \N__2577\ : std_logic;
signal \N__2574\ : std_logic;
signal \N__2571\ : std_logic;
signal \N__2568\ : std_logic;
signal \N__2563\ : std_logic;
signal \N__2560\ : std_logic;
signal \N__2557\ : std_logic;
signal \N__2554\ : std_logic;
signal \N__2553\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2547\ : std_logic;
signal \N__2544\ : std_logic;
signal \N__2539\ : std_logic;
signal \N__2538\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2521\ : std_logic;
signal \N__2518\ : std_logic;
signal \N__2515\ : std_logic;
signal \N__2512\ : std_logic;
signal \N__2509\ : std_logic;
signal \N__2506\ : std_logic;
signal \N__2503\ : std_logic;
signal \N__2500\ : std_logic;
signal \N__2497\ : std_logic;
signal \N__2496\ : std_logic;
signal \N__2493\ : std_logic;
signal \N__2490\ : std_logic;
signal \N__2489\ : std_logic;
signal \N__2488\ : std_logic;
signal \N__2485\ : std_logic;
signal \N__2484\ : std_logic;
signal \N__2481\ : std_logic;
signal \N__2480\ : std_logic;
signal \N__2477\ : std_logic;
signal \N__2474\ : std_logic;
signal \N__2471\ : std_logic;
signal \N__2470\ : std_logic;
signal \N__2469\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2463\ : std_logic;
signal \N__2458\ : std_logic;
signal \N__2455\ : std_logic;
signal \N__2452\ : std_logic;
signal \N__2447\ : std_logic;
signal \N__2444\ : std_logic;
signal \N__2431\ : std_logic;
signal \N__2428\ : std_logic;
signal \N__2427\ : std_logic;
signal \N__2426\ : std_logic;
signal \N__2425\ : std_logic;
signal \N__2422\ : std_logic;
signal \N__2421\ : std_logic;
signal \N__2420\ : std_logic;
signal \N__2419\ : std_logic;
signal \N__2418\ : std_logic;
signal \N__2417\ : std_logic;
signal \N__2414\ : std_logic;
signal \N__2409\ : std_logic;
signal \N__2406\ : std_logic;
signal \N__2403\ : std_logic;
signal \N__2400\ : std_logic;
signal \N__2397\ : std_logic;
signal \N__2392\ : std_logic;
signal \N__2389\ : std_logic;
signal \N__2374\ : std_logic;
signal \N__2371\ : std_logic;
signal \N__2370\ : std_logic;
signal \N__2369\ : std_logic;
signal \N__2368\ : std_logic;
signal \N__2367\ : std_logic;
signal \N__2366\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2362\ : std_logic;
signal \N__2361\ : std_logic;
signal \N__2358\ : std_logic;
signal \N__2355\ : std_logic;
signal \N__2352\ : std_logic;
signal \N__2347\ : std_logic;
signal \N__2344\ : std_logic;
signal \N__2339\ : std_logic;
signal \N__2336\ : std_logic;
signal \N__2323\ : std_logic;
signal \N__2322\ : std_logic;
signal \N__2319\ : std_logic;
signal \N__2318\ : std_logic;
signal \N__2315\ : std_logic;
signal \N__2314\ : std_logic;
signal \N__2313\ : std_logic;
signal \N__2312\ : std_logic;
signal \N__2309\ : std_logic;
signal \N__2306\ : std_logic;
signal \N__2305\ : std_logic;
signal \N__2304\ : std_logic;
signal \N__2301\ : std_logic;
signal \N__2298\ : std_logic;
signal \N__2293\ : std_logic;
signal \N__2290\ : std_logic;
signal \N__2287\ : std_logic;
signal \N__2284\ : std_logic;
signal \N__2281\ : std_logic;
signal \N__2266\ : std_logic;
signal \N__2263\ : std_logic;
signal \N__2260\ : std_logic;
signal \N__2257\ : std_logic;
signal \N__2254\ : std_logic;
signal \N__2251\ : std_logic;
signal \N__2248\ : std_logic;
signal \N__2245\ : std_logic;
signal \N__2242\ : std_logic;
signal \N__2239\ : std_logic;
signal \N__2236\ : std_logic;
signal \N__2233\ : std_logic;
signal \N__2230\ : std_logic;
signal \N__2227\ : std_logic;
signal \N__2226\ : std_logic;
signal \N__2225\ : std_logic;
signal \N__2222\ : std_logic;
signal \N__2221\ : std_logic;
signal \N__2220\ : std_logic;
signal \N__2217\ : std_logic;
signal \N__2210\ : std_logic;
signal \N__2209\ : std_logic;
signal \N__2204\ : std_logic;
signal \N__2203\ : std_logic;
signal \N__2202\ : std_logic;
signal \N__2201\ : std_logic;
signal \N__2200\ : std_logic;
signal \N__2199\ : std_logic;
signal \N__2198\ : std_logic;
signal \N__2197\ : std_logic;
signal \N__2194\ : std_logic;
signal \N__2191\ : std_logic;
signal \N__2188\ : std_logic;
signal \N__2185\ : std_logic;
signal \N__2182\ : std_logic;
signal \N__2179\ : std_logic;
signal \N__2176\ : std_logic;
signal \N__2173\ : std_logic;
signal \N__2170\ : std_logic;
signal \N__2167\ : std_logic;
signal \N__2164\ : std_logic;
signal \N__2161\ : std_logic;
signal \N__2158\ : std_logic;
signal \N__2151\ : std_logic;
signal \N__2142\ : std_logic;
signal \N__2131\ : std_logic;
signal \N__2128\ : std_logic;
signal \N__2125\ : std_logic;
signal \N__2122\ : std_logic;
signal \N__2119\ : std_logic;
signal \N__2116\ : std_logic;
signal \N__2113\ : std_logic;
signal \N__2110\ : std_logic;
signal \N__2107\ : std_logic;
signal \N__2106\ : std_logic;
signal \N__2101\ : std_logic;
signal \N__2098\ : std_logic;
signal \N__2095\ : std_logic;
signal \N__2092\ : std_logic;
signal \N__2089\ : std_logic;
signal \N__2086\ : std_logic;
signal \N__2083\ : std_logic;
signal \N__2080\ : std_logic;
signal \N__2077\ : std_logic;
signal \N__2074\ : std_logic;
signal \N__2071\ : std_logic;
signal \N__2068\ : std_logic;
signal \N__2065\ : std_logic;
signal \N__2064\ : std_logic;
signal \N__2063\ : std_logic;
signal \N__2060\ : std_logic;
signal \N__2057\ : std_logic;
signal \N__2054\ : std_logic;
signal \N__2051\ : std_logic;
signal \N__2044\ : std_logic;
signal \N__2041\ : std_logic;
signal \N__2038\ : std_logic;
signal \N__2035\ : std_logic;
signal \N__2034\ : std_logic;
signal \N__2033\ : std_logic;
signal \N__2030\ : std_logic;
signal \N__2027\ : std_logic;
signal \N__2024\ : std_logic;
signal \N__2021\ : std_logic;
signal \N__2018\ : std_logic;
signal \N__2011\ : std_logic;
signal \N__2008\ : std_logic;
signal \N__2005\ : std_logic;
signal \N__2002\ : std_logic;
signal \N__1999\ : std_logic;
signal \N__1996\ : std_logic;
signal \N__1993\ : std_logic;
signal \N__1990\ : std_logic;
signal \N__1987\ : std_logic;
signal \N__1984\ : std_logic;
signal \N__1981\ : std_logic;
signal \N__1978\ : std_logic;
signal \N__1975\ : std_logic;
signal \N__1972\ : std_logic;
signal \N__1969\ : std_logic;
signal \N__1966\ : std_logic;
signal \N__1963\ : std_logic;
signal \N__1962\ : std_logic;
signal \N__1961\ : std_logic;
signal \N__1956\ : std_logic;
signal \N__1953\ : std_logic;
signal \N__1948\ : std_logic;
signal \N__1945\ : std_logic;
signal \N__1942\ : std_logic;
signal \N__1939\ : std_logic;
signal \N__1936\ : std_logic;
signal \N__1933\ : std_logic;
signal \N__1932\ : std_logic;
signal \N__1931\ : std_logic;
signal \N__1928\ : std_logic;
signal \N__1923\ : std_logic;
signal \N__1918\ : std_logic;
signal \N__1915\ : std_logic;
signal \N__1912\ : std_logic;
signal \N__1909\ : std_logic;
signal \N__1906\ : std_logic;
signal \N__1903\ : std_logic;
signal \N__1900\ : std_logic;
signal \N__1899\ : std_logic;
signal \N__1898\ : std_logic;
signal \N__1895\ : std_logic;
signal \N__1890\ : std_logic;
signal \N__1885\ : std_logic;
signal \N__1882\ : std_logic;
signal \N__1879\ : std_logic;
signal \N__1876\ : std_logic;
signal \N__1873\ : std_logic;
signal \N__1870\ : std_logic;
signal \N__1867\ : std_logic;
signal \N__1864\ : std_logic;
signal \N__1861\ : std_logic;
signal \N__1858\ : std_logic;
signal \N__1855\ : std_logic;
signal \N__1852\ : std_logic;
signal \N__1849\ : std_logic;
signal \N__1848\ : std_logic;
signal \N__1845\ : std_logic;
signal \N__1842\ : std_logic;
signal \N__1841\ : std_logic;
signal \N__1838\ : std_logic;
signal \N__1833\ : std_logic;
signal \N__1828\ : std_logic;
signal \N__1827\ : std_logic;
signal \N__1824\ : std_logic;
signal \N__1821\ : std_logic;
signal \N__1820\ : std_logic;
signal \N__1817\ : std_logic;
signal \N__1814\ : std_logic;
signal \N__1811\ : std_logic;
signal \N__1804\ : std_logic;
signal \N__1803\ : std_logic;
signal \N__1800\ : std_logic;
signal \N__1799\ : std_logic;
signal \N__1796\ : std_logic;
signal \N__1793\ : std_logic;
signal \N__1788\ : std_logic;
signal \N__1783\ : std_logic;
signal \N__1780\ : std_logic;
signal \N__1779\ : std_logic;
signal \N__1778\ : std_logic;
signal \N__1775\ : std_logic;
signal \N__1770\ : std_logic;
signal \N__1765\ : std_logic;
signal \N__1762\ : std_logic;
signal \N__1759\ : std_logic;
signal \N__1756\ : std_logic;
signal \N__1753\ : std_logic;
signal \N__1750\ : std_logic;
signal \N__1747\ : std_logic;
signal \N__1744\ : std_logic;
signal \N__1743\ : std_logic;
signal \N__1740\ : std_logic;
signal \N__1737\ : std_logic;
signal \N__1732\ : std_logic;
signal \N__1731\ : std_logic;
signal \N__1728\ : std_logic;
signal \N__1725\ : std_logic;
signal \N__1722\ : std_logic;
signal \N__1717\ : std_logic;
signal \N__1714\ : std_logic;
signal \N__1711\ : std_logic;
signal \N__1710\ : std_logic;
signal \N__1709\ : std_logic;
signal \N__1706\ : std_logic;
signal \N__1701\ : std_logic;
signal \N__1696\ : std_logic;
signal \N__1693\ : std_logic;
signal \N__1690\ : std_logic;
signal \N__1687\ : std_logic;
signal \N__1684\ : std_logic;
signal \N__1683\ : std_logic;
signal \N__1680\ : std_logic;
signal \N__1677\ : std_logic;
signal \N__1672\ : std_logic;
signal \N__1669\ : std_logic;
signal \N__1666\ : std_logic;
signal \N__1663\ : std_logic;
signal \N__1662\ : std_logic;
signal \N__1659\ : std_logic;
signal \N__1656\ : std_logic;
signal \N__1651\ : std_logic;
signal \N__1648\ : std_logic;
signal \N__1645\ : std_logic;
signal \N__1642\ : std_logic;
signal \N__1641\ : std_logic;
signal \N__1638\ : std_logic;
signal \N__1635\ : std_logic;
signal \N__1630\ : std_logic;
signal \N__1627\ : std_logic;
signal \N__1624\ : std_logic;
signal \N__1621\ : std_logic;
signal \N__1620\ : std_logic;
signal \N__1617\ : std_logic;
signal \N__1614\ : std_logic;
signal \N__1609\ : std_logic;
signal \N__1606\ : std_logic;
signal \N__1603\ : std_logic;
signal \N__1600\ : std_logic;
signal \N__1599\ : std_logic;
signal \N__1596\ : std_logic;
signal \N__1593\ : std_logic;
signal \N__1588\ : std_logic;
signal \N__1585\ : std_logic;
signal \N__1582\ : std_logic;
signal \N__1579\ : std_logic;
signal \N__1578\ : std_logic;
signal \N__1575\ : std_logic;
signal \N__1572\ : std_logic;
signal \N__1567\ : std_logic;
signal \N__1564\ : std_logic;
signal \N__1561\ : std_logic;
signal \N__1560\ : std_logic;
signal \N__1557\ : std_logic;
signal \N__1554\ : std_logic;
signal \N__1549\ : std_logic;
signal \N__1546\ : std_logic;
signal \N__1543\ : std_logic;
signal \N__1540\ : std_logic;
signal \N__1537\ : std_logic;
signal \N__1534\ : std_logic;
signal \N__1531\ : std_logic;
signal \N__1528\ : std_logic;
signal \N__1525\ : std_logic;
signal \N__1522\ : std_logic;
signal \N__1519\ : std_logic;
signal \N__1516\ : std_logic;
signal \N__1513\ : std_logic;
signal \N__1510\ : std_logic;
signal \N__1507\ : std_logic;
signal \N__1504\ : std_logic;
signal \N__1501\ : std_logic;
signal \N__1498\ : std_logic;
signal \N__1495\ : std_logic;
signal \N__1492\ : std_logic;
signal \N__1489\ : std_logic;
signal \N__1486\ : std_logic;
signal \N__1483\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \my_uart.recv_state_0_sqmuxa_1_cascade_\ : std_logic;
signal \my_uart.g0_2\ : std_logic;
signal \my_uart.g0_0_0_a3_0_0_cascade_\ : std_logic;
signal \my_uart.g0_0_0_a3_0_4\ : std_logic;
signal \my_uart.rx_bits_remaining_6_0_3\ : std_logic;
signal \my_uart.g0_0_0_a3_3_cascade_\ : std_logic;
signal \my_uart.N_4_cascade_\ : std_logic;
signal \my_uart.g0_0\ : std_logic;
signal \my_uart.g0_0_0_a3_4\ : std_logic;
signal \LED_o_c_0\ : std_logic;
signal \LED_o_c_7\ : std_logic;
signal \LED_o_c_6\ : std_logic;
signal \LED_o_c_3\ : std_logic;
signal \LED_o_c_2\ : std_logic;
signal \LED_o_c_1\ : std_logic;
signal \LED_o_c_5\ : std_logic;
signal \LED_o_c_4\ : std_logic;
signal \bfn_9_25_0_\ : std_logic;
signal \my_uart.rx_clk_divider_1_cry_0\ : std_logic;
signal \my_uart.rx_clk_divider_1_cry_1\ : std_logic;
signal \my_uart.rx_clk_divider_1_cry_2\ : std_logic;
signal \my_uart.rx_clk_divider_1_cry_3\ : std_logic;
signal \my_uart.rx_clk_divider_1_cry_4\ : std_logic;
signal \my_uart.rx_clk_divider_1_cry_5\ : std_logic;
signal \my_uart.rx_clk_divider_1_cry_6\ : std_logic;
signal \my_uart.rx_clk_divider_1_cry_7\ : std_logic;
signal \bfn_9_26_0_\ : std_logic;
signal \my_uart.rx_clk_divider_1_cry_8\ : std_logic;
signal \my_uart.rx_clk_divider_1_cry_9\ : std_logic;
signal \my_uart.rx_clk_dividerZ0Z_1\ : std_logic;
signal \my_uart.rx_clk_dividerZ0Z_10\ : std_logic;
signal \my_uart.rx_clk_divider_1_cry_0_THRU_CO\ : std_logic;
signal \my_uart.rx_clk_dividerZ1Z_1\ : std_logic;
signal \my_uart.rx_clk_divider_1_cry_7_THRU_CO\ : std_logic;
signal \my_uart.rx_clk_divider_1_cry_8_THRU_CO\ : std_logic;
signal \my_uart.rx_clk_divider_1_cry_1_THRU_CO\ : std_logic;
signal \my_uart.rx_clk_dividerZ0Z_2\ : std_logic;
signal \my_uart.rx_clk_divider_1_cry_2_THRU_CO\ : std_logic;
signal \my_uart.rx_clk_divider_1_cry_3_THRU_CO\ : std_logic;
signal \my_uart.rx_clk_divider_1_cry_5_THRU_CO\ : std_logic;
signal \my_uart.rx_clk_divider_1_cry_4_THRU_CO\ : std_logic;
signal \my_uart.rx_clk_dividerZ0Z_5\ : std_logic;
signal \my_uart.rx_clk_dividerZ0Z_4\ : std_logic;
signal \my_uart.rx_clk_dividerZ0Z_6\ : std_logic;
signal \my_uart.rx_clk_dividerZ0Z_3\ : std_logic;
signal \my_uart.rx_countdown_8_5_cascade_\ : std_logic;
signal \my_uart.rx_clk_dividerZ0Z_8\ : std_logic;
signal \my_uart.rx_countdown_RNO_5Z0Z_2\ : std_logic;
signal \my_uart.rx_countdown_RNO_6Z0Z_2_cascade_\ : std_logic;
signal \my_uart.rx_clk_divider_1_cry_6_THRU_CO\ : std_logic;
signal \my_uart.rx_clk_dividerZ0Z_7\ : std_logic;
signal \my_uart.rx_data_0_sqmuxa\ : std_logic;
signal \my_uart.N_6_cascade_\ : std_logic;
signal \my_uart.un1_rx_clk_divider_a_0\ : std_logic;
signal \my_uart.rx_clk_dividerZ0Z_9\ : std_logic;
signal \my_uart.un1_rx_clk_divider_a_6\ : std_logic;
signal \my_uart.un1_rx_clk_divider_a_7\ : std_logic;
signal \my_uart.un1_rx_clk_divider_a_cascade_\ : std_logic;
signal \my_uart.N_5\ : std_logic;
signal \my_uart.g0_0_0_a3_0_3\ : std_logic;
signal \my_uart.g0_6_a5_1_5_cascade_\ : std_logic;
signal \my_uart.g0_6_a5_1_4\ : std_logic;
signal \my_uart.rx_countdown_3_4\ : std_logic;
signal \my_uart.rx_countdown_3_4_cascade_\ : std_logic;
signal \my_uart.rx_countdown_RNO_4Z0Z_2\ : std_logic;
signal \my_uart.N_13\ : std_logic;
signal \my_uart.rx_countdown_3_3\ : std_logic;
signal \my_uart.G_14_0_a3_0_1\ : std_logic;
signal \my_uart.g0_6_0_0\ : std_logic;
signal \my_uart.g0_4_a3_0_3\ : std_logic;
signal \my_uart.rx_countdown20_cascade_\ : std_logic;
signal \my_uart.un1_recv_state_6\ : std_logic;
signal \my_uart.g0_4_a3_3_cascade_\ : std_logic;
signal \my_uart.g0_4_a3_4\ : std_logic;
signal \my_uart.recv_state_0_sqmuxa_1_0\ : std_logic;
signal \my_uart.g0_4_a3_0_2\ : std_logic;
signal \my_uart.g0_6_a5_1_0\ : std_logic;
signal \bfn_11_26_0_\ : std_logic;
signal \my_uart.rx_countdown_3_cry_0_s1\ : std_logic;
signal \my_uart.rx_countdown_3_cry_1_s1\ : std_logic;
signal \my_uart.rx_countdown_3_cry_2_s1\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \my_uart.rx_countdown_3_cry_3_s1\ : std_logic;
signal \my_uart.rx_countdown_3_cry_4_s1\ : std_logic;
signal \my_uart.un1_recv_state_8\ : std_logic;
signal \my_uart.g0_0_0_a3_3_0\ : std_logic;
signal \my_uart.N_8_0_cascade_\ : std_logic;
signal \my_uart.N_18_mux\ : std_logic;
signal \my_uart.rx_countdownZ0Z_4\ : std_logic;
signal \my_uart.rx_countdownZ1Z_1\ : std_logic;
signal \my_uart.rx_countdownZ1Z_2\ : std_logic;
signal \my_uart.rx_countdownZ1Z_3\ : std_logic;
signal \my_uart.m10_e_1_cascade_\ : std_logic;
signal \my_uart.rx_countdownZ0Z_5\ : std_logic;
signal \my_uart.N_22_mux\ : std_logic;
signal \my_uart.N_23_mux_cascade_\ : std_logic;
signal \my_uart.m7_0_0\ : std_logic;
signal \my_uart.g0_6_0_1\ : std_logic;
signal \my_uart.un1_rx_clk_divider28_i_cascade_\ : std_logic;
signal \my_uart.rx_clk_divider_0_sqmuxa\ : std_logic;
signal \my_uart.m6_0_18_0\ : std_logic;
signal \my_uart.rx_bits_remainingZ0Z_3\ : std_logic;
signal \my_uart.rx_bits_remainingZ0Z_1\ : std_logic;
signal \my_uart.rx_bits_remainingZ0Z_0\ : std_logic;
signal \my_uart.CO1_i\ : std_logic;
signal \my_uart.CO1_i_cascade_\ : std_logic;
signal \my_uart.rx_bits_remainingZ0Z_2\ : std_logic;
signal \my_uart.un1_rx_data_0_sqmuxa_i_i\ : std_logic;
signal \CLK_i_c_g\ : std_logic;
signal \my_uart.m15_e_0_cascade_\ : std_logic;
signal \my_uart.m15_e_3_cascade_\ : std_logic;
signal \my_uart.N_28_mux\ : std_logic;
signal \my_uart.N_19_mux_0\ : std_logic;
signal \my_uart.m10_e_3\ : std_logic;
signal \my_uart.N_19_mux_0_cascade_\ : std_logic;
signal \my_uart.un1_rx_clk_divider_a\ : std_logic;
signal \my_uart.N_27_mux\ : std_logic;
signal \RS232_RX_i_c\ : std_logic;
signal \N_20_mux\ : std_logic;
signal \my_uart.N_11\ : std_logic;
signal \my_uart.rx_countdown_3_s1_3\ : std_logic;
signal \my_uart.g0_6_a5_0_5\ : std_logic;
signal \my_uart.rx_countdownZ0Z_3\ : std_logic;
signal \my_uart.N_19_mux\ : std_logic;
signal \my_uart.m6_0_18_a4_1_2\ : std_logic;
signal my_uart_recv_state_2 : std_logic;
signal \my_uart.N_217\ : std_logic;
signal \N_18_i\ : std_logic;
signal \my_uart.rx_countdown_3_s1_1\ : std_logic;
signal my_uart_recv_state_0 : std_logic;
signal \my_uart.rx_countdown_3_s1_2\ : std_logic;
signal \my_uart.g0_6_a5_0_4\ : std_logic;
signal \my_uart.rx_countdown_3_s1_4\ : std_logic;
signal \my_uart.rx_countdown_3_s1_5\ : std_logic;
signal \my_uart.g0_6_a5_0_3\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK_i_wire\ : std_logic;
signal \LED_o_wire\ : std_logic_vector(7 downto 0);
signal \RS232_RX_i_wire\ : std_logic;

begin
    \CLK_i_wire\ <= CLK_i;
    LED_o <= \LED_o_wire\;
    \RS232_RX_i_wire\ <= RS232_RX_i;

    \CLK_i_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__3941\,
            GLOBALBUFFEROUTPUT => \CLK_i_c_g\
        );

    \CLK_i_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3943\,
            DIN => \N__3942\,
            DOUT => \N__3941\,
            PACKAGEPIN => \CLK_i_wire\
        );

    \CLK_i_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3943\,
            PADOUT => \N__3942\,
            PADIN => \N__3941\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED_o_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3932\,
            DIN => \N__3931\,
            DOUT => \N__3930\,
            PACKAGEPIN => \LED_o_wire\(0)
        );

    \LED_o_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3932\,
            PADOUT => \N__3931\,
            PADIN => \N__3930\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1513\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED_o_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3923\,
            DIN => \N__3922\,
            DOUT => \N__3921\,
            PACKAGEPIN => \LED_o_wire\(5)
        );

    \LED_o_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3923\,
            PADOUT => \N__3922\,
            PADIN => \N__3921\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1588\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED_o_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3914\,
            DIN => \N__3913\,
            DOUT => \N__3912\,
            PACKAGEPIN => \LED_o_wire\(1)
        );

    \LED_o_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3914\,
            PADOUT => \N__3913\,
            PADIN => \N__3912\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1609\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED_o_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3905\,
            DIN => \N__3904\,
            DOUT => \N__3903\,
            PACKAGEPIN => \LED_o_wire\(6)
        );

    \LED_o_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3905\,
            PADOUT => \N__3904\,
            PADIN => \N__3903\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1672\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED_o_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3896\,
            DIN => \N__3895\,
            DOUT => \N__3894\,
            PACKAGEPIN => \LED_o_wire\(2)
        );

    \LED_o_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3896\,
            PADOUT => \N__3895\,
            PADIN => \N__3894\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1630\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RS232_RX_i_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3887\,
            DIN => \N__3886\,
            DOUT => \N__3885\,
            PACKAGEPIN => \RS232_RX_i_wire\
        );

    \RS232_RX_i_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3887\,
            PADOUT => \N__3886\,
            PADIN => \N__3885\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RS232_RX_i_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED_o_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3878\,
            DIN => \N__3877\,
            DOUT => \N__3876\,
            PACKAGEPIN => \LED_o_wire\(7)
        );

    \LED_o_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3878\,
            PADOUT => \N__3877\,
            PADIN => \N__3876\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1696\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED_o_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3869\,
            DIN => \N__3868\,
            DOUT => \N__3867\,
            PACKAGEPIN => \LED_o_wire\(3)
        );

    \LED_o_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3869\,
            PADOUT => \N__3868\,
            PADIN => \N__3867\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1651\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED_o_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3860\,
            DIN => \N__3859\,
            DOUT => \N__3858\,
            PACKAGEPIN => \LED_o_wire\(4)
        );

    \LED_o_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3860\,
            PADOUT => \N__3859\,
            PADIN => \N__3858\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1567\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__913\ : CascadeMux
    port map (
            O => \N__3841\,
            I => \N__3838\
        );

    \I__912\ : InMux
    port map (
            O => \N__3838\,
            I => \N__3835\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__3835\,
            I => \N__3825\
        );

    \I__910\ : InMux
    port map (
            O => \N__3834\,
            I => \N__3822\
        );

    \I__909\ : InMux
    port map (
            O => \N__3833\,
            I => \N__3819\
        );

    \I__908\ : CascadeMux
    port map (
            O => \N__3832\,
            I => \N__3816\
        );

    \I__907\ : CascadeMux
    port map (
            O => \N__3831\,
            I => \N__3813\
        );

    \I__906\ : CascadeMux
    port map (
            O => \N__3830\,
            I => \N__3810\
        );

    \I__905\ : CascadeMux
    port map (
            O => \N__3829\,
            I => \N__3807\
        );

    \I__904\ : CascadeMux
    port map (
            O => \N__3828\,
            I => \N__3803\
        );

    \I__903\ : Span4Mux_v
    port map (
            O => \N__3825\,
            I => \N__3798\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__3822\,
            I => \N__3798\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__3819\,
            I => \N__3795\
        );

    \I__900\ : InMux
    port map (
            O => \N__3816\,
            I => \N__3790\
        );

    \I__899\ : InMux
    port map (
            O => \N__3813\,
            I => \N__3790\
        );

    \I__898\ : InMux
    port map (
            O => \N__3810\,
            I => \N__3785\
        );

    \I__897\ : InMux
    port map (
            O => \N__3807\,
            I => \N__3785\
        );

    \I__896\ : InMux
    port map (
            O => \N__3806\,
            I => \N__3782\
        );

    \I__895\ : InMux
    port map (
            O => \N__3803\,
            I => \N__3779\
        );

    \I__894\ : Span4Mux_v
    port map (
            O => \N__3798\,
            I => \N__3776\
        );

    \I__893\ : Span4Mux_v
    port map (
            O => \N__3795\,
            I => \N__3773\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__3790\,
            I => \N__3768\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__3785\,
            I => \N__3768\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__3782\,
            I => \N__3765\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__3779\,
            I => \N__3762\
        );

    \I__888\ : Span4Mux_h
    port map (
            O => \N__3776\,
            I => \N__3755\
        );

    \I__887\ : Span4Mux_s3_v
    port map (
            O => \N__3773\,
            I => \N__3755\
        );

    \I__886\ : Span4Mux_v
    port map (
            O => \N__3768\,
            I => \N__3755\
        );

    \I__885\ : Sp12to4
    port map (
            O => \N__3765\,
            I => \N__3752\
        );

    \I__884\ : Span12Mux_v
    port map (
            O => \N__3762\,
            I => \N__3747\
        );

    \I__883\ : Sp12to4
    port map (
            O => \N__3755\,
            I => \N__3747\
        );

    \I__882\ : Span12Mux_h
    port map (
            O => \N__3752\,
            I => \N__3744\
        );

    \I__881\ : Span12Mux_h
    port map (
            O => \N__3747\,
            I => \N__3741\
        );

    \I__880\ : Odrv12
    port map (
            O => \N__3744\,
            I => \RS232_RX_i_c\
        );

    \I__879\ : Odrv12
    port map (
            O => \N__3741\,
            I => \RS232_RX_i_c\
        );

    \I__878\ : InMux
    port map (
            O => \N__3736\,
            I => \N__3730\
        );

    \I__877\ : InMux
    port map (
            O => \N__3735\,
            I => \N__3730\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__3730\,
            I => \N_20_mux\
        );

    \I__875\ : InMux
    port map (
            O => \N__3727\,
            I => \N__3724\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__3724\,
            I => \N__3721\
        );

    \I__873\ : Odrv4
    port map (
            O => \N__3721\,
            I => \my_uart.N_11\
        );

    \I__872\ : InMux
    port map (
            O => \N__3718\,
            I => \N__3711\
        );

    \I__871\ : InMux
    port map (
            O => \N__3717\,
            I => \N__3706\
        );

    \I__870\ : InMux
    port map (
            O => \N__3716\,
            I => \N__3703\
        );

    \I__869\ : InMux
    port map (
            O => \N__3715\,
            I => \N__3700\
        );

    \I__868\ : InMux
    port map (
            O => \N__3714\,
            I => \N__3697\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__3711\,
            I => \N__3694\
        );

    \I__866\ : InMux
    port map (
            O => \N__3710\,
            I => \N__3691\
        );

    \I__865\ : InMux
    port map (
            O => \N__3709\,
            I => \N__3688\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__3706\,
            I => \my_uart.rx_countdown_3_s1_3\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__3703\,
            I => \my_uart.rx_countdown_3_s1_3\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__3700\,
            I => \my_uart.rx_countdown_3_s1_3\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__3697\,
            I => \my_uart.rx_countdown_3_s1_3\
        );

    \I__860\ : Odrv12
    port map (
            O => \N__3694\,
            I => \my_uart.rx_countdown_3_s1_3\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__3691\,
            I => \my_uart.rx_countdown_3_s1_3\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__3688\,
            I => \my_uart.rx_countdown_3_s1_3\
        );

    \I__857\ : InMux
    port map (
            O => \N__3673\,
            I => \N__3670\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__3670\,
            I => \my_uart.g0_6_a5_0_5\
        );

    \I__855\ : InMux
    port map (
            O => \N__3667\,
            I => \N__3663\
        );

    \I__854\ : InMux
    port map (
            O => \N__3666\,
            I => \N__3651\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__3663\,
            I => \N__3648\
        );

    \I__852\ : CascadeMux
    port map (
            O => \N__3662\,
            I => \N__3642\
        );

    \I__851\ : InMux
    port map (
            O => \N__3661\,
            I => \N__3639\
        );

    \I__850\ : InMux
    port map (
            O => \N__3660\,
            I => \N__3634\
        );

    \I__849\ : InMux
    port map (
            O => \N__3659\,
            I => \N__3634\
        );

    \I__848\ : InMux
    port map (
            O => \N__3658\,
            I => \N__3629\
        );

    \I__847\ : InMux
    port map (
            O => \N__3657\,
            I => \N__3629\
        );

    \I__846\ : InMux
    port map (
            O => \N__3656\,
            I => \N__3624\
        );

    \I__845\ : InMux
    port map (
            O => \N__3655\,
            I => \N__3624\
        );

    \I__844\ : InMux
    port map (
            O => \N__3654\,
            I => \N__3621\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__3651\,
            I => \N__3618\
        );

    \I__842\ : Span4Mux_h
    port map (
            O => \N__3648\,
            I => \N__3615\
        );

    \I__841\ : InMux
    port map (
            O => \N__3647\,
            I => \N__3612\
        );

    \I__840\ : InMux
    port map (
            O => \N__3646\,
            I => \N__3605\
        );

    \I__839\ : InMux
    port map (
            O => \N__3645\,
            I => \N__3605\
        );

    \I__838\ : InMux
    port map (
            O => \N__3642\,
            I => \N__3605\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__3639\,
            I => \my_uart.rx_countdownZ0Z_3\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__3634\,
            I => \my_uart.rx_countdownZ0Z_3\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__3629\,
            I => \my_uart.rx_countdownZ0Z_3\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__3624\,
            I => \my_uart.rx_countdownZ0Z_3\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__3621\,
            I => \my_uart.rx_countdownZ0Z_3\
        );

    \I__832\ : Odrv12
    port map (
            O => \N__3618\,
            I => \my_uart.rx_countdownZ0Z_3\
        );

    \I__831\ : Odrv4
    port map (
            O => \N__3615\,
            I => \my_uart.rx_countdownZ0Z_3\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__3612\,
            I => \my_uart.rx_countdownZ0Z_3\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__3605\,
            I => \my_uart.rx_countdownZ0Z_3\
        );

    \I__828\ : InMux
    port map (
            O => \N__3586\,
            I => \N__3583\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__3583\,
            I => \my_uart.N_19_mux\
        );

    \I__826\ : InMux
    port map (
            O => \N__3580\,
            I => \N__3577\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__3577\,
            I => \N__3574\
        );

    \I__824\ : Span4Mux_h
    port map (
            O => \N__3574\,
            I => \N__3571\
        );

    \I__823\ : Odrv4
    port map (
            O => \N__3571\,
            I => \my_uart.m6_0_18_a4_1_2\
        );

    \I__822\ : InMux
    port map (
            O => \N__3568\,
            I => \N__3564\
        );

    \I__821\ : InMux
    port map (
            O => \N__3567\,
            I => \N__3561\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__3564\,
            I => \N__3549\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__3561\,
            I => \N__3549\
        );

    \I__818\ : InMux
    port map (
            O => \N__3560\,
            I => \N__3544\
        );

    \I__817\ : InMux
    port map (
            O => \N__3559\,
            I => \N__3544\
        );

    \I__816\ : CascadeMux
    port map (
            O => \N__3558\,
            I => \N__3541\
        );

    \I__815\ : CascadeMux
    port map (
            O => \N__3557\,
            I => \N__3534\
        );

    \I__814\ : CascadeMux
    port map (
            O => \N__3556\,
            I => \N__3527\
        );

    \I__813\ : InMux
    port map (
            O => \N__3555\,
            I => \N__3522\
        );

    \I__812\ : InMux
    port map (
            O => \N__3554\,
            I => \N__3522\
        );

    \I__811\ : Span4Mux_v
    port map (
            O => \N__3549\,
            I => \N__3517\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__3544\,
            I => \N__3517\
        );

    \I__809\ : InMux
    port map (
            O => \N__3541\,
            I => \N__3513\
        );

    \I__808\ : InMux
    port map (
            O => \N__3540\,
            I => \N__3506\
        );

    \I__807\ : InMux
    port map (
            O => \N__3539\,
            I => \N__3506\
        );

    \I__806\ : InMux
    port map (
            O => \N__3538\,
            I => \N__3506\
        );

    \I__805\ : InMux
    port map (
            O => \N__3537\,
            I => \N__3501\
        );

    \I__804\ : InMux
    port map (
            O => \N__3534\,
            I => \N__3501\
        );

    \I__803\ : InMux
    port map (
            O => \N__3533\,
            I => \N__3494\
        );

    \I__802\ : InMux
    port map (
            O => \N__3532\,
            I => \N__3494\
        );

    \I__801\ : InMux
    port map (
            O => \N__3531\,
            I => \N__3494\
        );

    \I__800\ : InMux
    port map (
            O => \N__3530\,
            I => \N__3489\
        );

    \I__799\ : InMux
    port map (
            O => \N__3527\,
            I => \N__3489\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__3522\,
            I => \N__3484\
        );

    \I__797\ : Span4Mux_h
    port map (
            O => \N__3517\,
            I => \N__3484\
        );

    \I__796\ : InMux
    port map (
            O => \N__3516\,
            I => \N__3481\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__3513\,
            I => my_uart_recv_state_2
        );

    \I__794\ : LocalMux
    port map (
            O => \N__3506\,
            I => my_uart_recv_state_2
        );

    \I__793\ : LocalMux
    port map (
            O => \N__3501\,
            I => my_uart_recv_state_2
        );

    \I__792\ : LocalMux
    port map (
            O => \N__3494\,
            I => my_uart_recv_state_2
        );

    \I__791\ : LocalMux
    port map (
            O => \N__3489\,
            I => my_uart_recv_state_2
        );

    \I__790\ : Odrv4
    port map (
            O => \N__3484\,
            I => my_uart_recv_state_2
        );

    \I__789\ : LocalMux
    port map (
            O => \N__3481\,
            I => my_uart_recv_state_2
        );

    \I__788\ : InMux
    port map (
            O => \N__3466\,
            I => \N__3463\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__3463\,
            I => \my_uart.N_217\
        );

    \I__786\ : InMux
    port map (
            O => \N__3460\,
            I => \N__3455\
        );

    \I__785\ : CascadeMux
    port map (
            O => \N__3459\,
            I => \N__3451\
        );

    \I__784\ : CascadeMux
    port map (
            O => \N__3458\,
            I => \N__3448\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__3455\,
            I => \N__3444\
        );

    \I__782\ : InMux
    port map (
            O => \N__3454\,
            I => \N__3441\
        );

    \I__781\ : InMux
    port map (
            O => \N__3451\,
            I => \N__3429\
        );

    \I__780\ : InMux
    port map (
            O => \N__3448\,
            I => \N__3429\
        );

    \I__779\ : InMux
    port map (
            O => \N__3447\,
            I => \N__3429\
        );

    \I__778\ : Span4Mux_v
    port map (
            O => \N__3444\,
            I => \N__3424\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__3441\,
            I => \N__3424\
        );

    \I__776\ : InMux
    port map (
            O => \N__3440\,
            I => \N__3416\
        );

    \I__775\ : InMux
    port map (
            O => \N__3439\,
            I => \N__3413\
        );

    \I__774\ : InMux
    port map (
            O => \N__3438\,
            I => \N__3408\
        );

    \I__773\ : InMux
    port map (
            O => \N__3437\,
            I => \N__3408\
        );

    \I__772\ : InMux
    port map (
            O => \N__3436\,
            I => \N__3405\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__3429\,
            I => \N__3402\
        );

    \I__770\ : Span4Mux_h
    port map (
            O => \N__3424\,
            I => \N__3399\
        );

    \I__769\ : InMux
    port map (
            O => \N__3423\,
            I => \N__3394\
        );

    \I__768\ : InMux
    port map (
            O => \N__3422\,
            I => \N__3394\
        );

    \I__767\ : InMux
    port map (
            O => \N__3421\,
            I => \N__3391\
        );

    \I__766\ : InMux
    port map (
            O => \N__3420\,
            I => \N__3386\
        );

    \I__765\ : InMux
    port map (
            O => \N__3419\,
            I => \N__3386\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__3416\,
            I => \N_18_i\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__3413\,
            I => \N_18_i\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__3408\,
            I => \N_18_i\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__3405\,
            I => \N_18_i\
        );

    \I__760\ : Odrv4
    port map (
            O => \N__3402\,
            I => \N_18_i\
        );

    \I__759\ : Odrv4
    port map (
            O => \N__3399\,
            I => \N_18_i\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__3394\,
            I => \N_18_i\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__3391\,
            I => \N_18_i\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__3386\,
            I => \N_18_i\
        );

    \I__755\ : CascadeMux
    port map (
            O => \N__3367\,
            I => \N__3364\
        );

    \I__754\ : InMux
    port map (
            O => \N__3364\,
            I => \N__3355\
        );

    \I__753\ : CascadeMux
    port map (
            O => \N__3363\,
            I => \N__3351\
        );

    \I__752\ : CascadeMux
    port map (
            O => \N__3362\,
            I => \N__3348\
        );

    \I__751\ : InMux
    port map (
            O => \N__3361\,
            I => \N__3345\
        );

    \I__750\ : InMux
    port map (
            O => \N__3360\,
            I => \N__3340\
        );

    \I__749\ : InMux
    port map (
            O => \N__3359\,
            I => \N__3340\
        );

    \I__748\ : InMux
    port map (
            O => \N__3358\,
            I => \N__3337\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__3355\,
            I => \N__3334\
        );

    \I__746\ : InMux
    port map (
            O => \N__3354\,
            I => \N__3331\
        );

    \I__745\ : InMux
    port map (
            O => \N__3351\,
            I => \N__3328\
        );

    \I__744\ : InMux
    port map (
            O => \N__3348\,
            I => \N__3325\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__3345\,
            I => \my_uart.rx_countdown_3_s1_1\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__3340\,
            I => \my_uart.rx_countdown_3_s1_1\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__3337\,
            I => \my_uart.rx_countdown_3_s1_1\
        );

    \I__740\ : Odrv12
    port map (
            O => \N__3334\,
            I => \my_uart.rx_countdown_3_s1_1\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__3331\,
            I => \my_uart.rx_countdown_3_s1_1\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__3328\,
            I => \my_uart.rx_countdown_3_s1_1\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__3325\,
            I => \my_uart.rx_countdown_3_s1_1\
        );

    \I__736\ : InMux
    port map (
            O => \N__3310\,
            I => \N__3307\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__3307\,
            I => \N__3294\
        );

    \I__734\ : InMux
    port map (
            O => \N__3306\,
            I => \N__3289\
        );

    \I__733\ : InMux
    port map (
            O => \N__3305\,
            I => \N__3289\
        );

    \I__732\ : CascadeMux
    port map (
            O => \N__3304\,
            I => \N__3283\
        );

    \I__731\ : InMux
    port map (
            O => \N__3303\,
            I => \N__3275\
        );

    \I__730\ : InMux
    port map (
            O => \N__3302\,
            I => \N__3275\
        );

    \I__729\ : InMux
    port map (
            O => \N__3301\,
            I => \N__3275\
        );

    \I__728\ : CascadeMux
    port map (
            O => \N__3300\,
            I => \N__3268\
        );

    \I__727\ : InMux
    port map (
            O => \N__3299\,
            I => \N__3261\
        );

    \I__726\ : InMux
    port map (
            O => \N__3298\,
            I => \N__3261\
        );

    \I__725\ : InMux
    port map (
            O => \N__3297\,
            I => \N__3261\
        );

    \I__724\ : Span4Mux_v
    port map (
            O => \N__3294\,
            I => \N__3256\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__3289\,
            I => \N__3256\
        );

    \I__722\ : InMux
    port map (
            O => \N__3288\,
            I => \N__3249\
        );

    \I__721\ : InMux
    port map (
            O => \N__3287\,
            I => \N__3249\
        );

    \I__720\ : InMux
    port map (
            O => \N__3286\,
            I => \N__3249\
        );

    \I__719\ : InMux
    port map (
            O => \N__3283\,
            I => \N__3246\
        );

    \I__718\ : InMux
    port map (
            O => \N__3282\,
            I => \N__3241\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__3275\,
            I => \N__3238\
        );

    \I__716\ : InMux
    port map (
            O => \N__3274\,
            I => \N__3231\
        );

    \I__715\ : InMux
    port map (
            O => \N__3273\,
            I => \N__3231\
        );

    \I__714\ : InMux
    port map (
            O => \N__3272\,
            I => \N__3231\
        );

    \I__713\ : InMux
    port map (
            O => \N__3271\,
            I => \N__3226\
        );

    \I__712\ : InMux
    port map (
            O => \N__3268\,
            I => \N__3226\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__3261\,
            I => \N__3223\
        );

    \I__710\ : Span4Mux_h
    port map (
            O => \N__3256\,
            I => \N__3220\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__3249\,
            I => \N__3217\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__3246\,
            I => \N__3214\
        );

    \I__707\ : InMux
    port map (
            O => \N__3245\,
            I => \N__3209\
        );

    \I__706\ : InMux
    port map (
            O => \N__3244\,
            I => \N__3209\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__3241\,
            I => my_uart_recv_state_0
        );

    \I__704\ : Odrv4
    port map (
            O => \N__3238\,
            I => my_uart_recv_state_0
        );

    \I__703\ : LocalMux
    port map (
            O => \N__3231\,
            I => my_uart_recv_state_0
        );

    \I__702\ : LocalMux
    port map (
            O => \N__3226\,
            I => my_uart_recv_state_0
        );

    \I__701\ : Odrv4
    port map (
            O => \N__3223\,
            I => my_uart_recv_state_0
        );

    \I__700\ : Odrv4
    port map (
            O => \N__3220\,
            I => my_uart_recv_state_0
        );

    \I__699\ : Odrv4
    port map (
            O => \N__3217\,
            I => my_uart_recv_state_0
        );

    \I__698\ : Odrv4
    port map (
            O => \N__3214\,
            I => my_uart_recv_state_0
        );

    \I__697\ : LocalMux
    port map (
            O => \N__3209\,
            I => my_uart_recv_state_0
        );

    \I__696\ : InMux
    port map (
            O => \N__3190\,
            I => \N__3182\
        );

    \I__695\ : InMux
    port map (
            O => \N__3189\,
            I => \N__3179\
        );

    \I__694\ : InMux
    port map (
            O => \N__3188\,
            I => \N__3175\
        );

    \I__693\ : InMux
    port map (
            O => \N__3187\,
            I => \N__3172\
        );

    \I__692\ : InMux
    port map (
            O => \N__3186\,
            I => \N__3169\
        );

    \I__691\ : InMux
    port map (
            O => \N__3185\,
            I => \N__3166\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__3182\,
            I => \N__3163\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__3179\,
            I => \N__3160\
        );

    \I__688\ : InMux
    port map (
            O => \N__3178\,
            I => \N__3157\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__3175\,
            I => \my_uart.rx_countdown_3_s1_2\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__3172\,
            I => \my_uart.rx_countdown_3_s1_2\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__3169\,
            I => \my_uart.rx_countdown_3_s1_2\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__3166\,
            I => \my_uart.rx_countdown_3_s1_2\
        );

    \I__683\ : Odrv12
    port map (
            O => \N__3163\,
            I => \my_uart.rx_countdown_3_s1_2\
        );

    \I__682\ : Odrv12
    port map (
            O => \N__3160\,
            I => \my_uart.rx_countdown_3_s1_2\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__3157\,
            I => \my_uart.rx_countdown_3_s1_2\
        );

    \I__680\ : CascadeMux
    port map (
            O => \N__3142\,
            I => \N__3139\
        );

    \I__679\ : InMux
    port map (
            O => \N__3139\,
            I => \N__3136\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__3136\,
            I => \my_uart.g0_6_a5_0_4\
        );

    \I__677\ : InMux
    port map (
            O => \N__3133\,
            I => \N__3125\
        );

    \I__676\ : InMux
    port map (
            O => \N__3132\,
            I => \N__3125\
        );

    \I__675\ : InMux
    port map (
            O => \N__3131\,
            I => \N__3119\
        );

    \I__674\ : InMux
    port map (
            O => \N__3130\,
            I => \N__3116\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__3125\,
            I => \N__3113\
        );

    \I__672\ : InMux
    port map (
            O => \N__3124\,
            I => \N__3110\
        );

    \I__671\ : InMux
    port map (
            O => \N__3123\,
            I => \N__3107\
        );

    \I__670\ : InMux
    port map (
            O => \N__3122\,
            I => \N__3104\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__3119\,
            I => \my_uart.rx_countdown_3_s1_4\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__3116\,
            I => \my_uart.rx_countdown_3_s1_4\
        );

    \I__667\ : Odrv12
    port map (
            O => \N__3113\,
            I => \my_uart.rx_countdown_3_s1_4\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__3110\,
            I => \my_uart.rx_countdown_3_s1_4\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3107\,
            I => \my_uart.rx_countdown_3_s1_4\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__3104\,
            I => \my_uart.rx_countdown_3_s1_4\
        );

    \I__663\ : InMux
    port map (
            O => \N__3091\,
            I => \N__3083\
        );

    \I__662\ : InMux
    port map (
            O => \N__3090\,
            I => \N__3083\
        );

    \I__661\ : InMux
    port map (
            O => \N__3089\,
            I => \N__3076\
        );

    \I__660\ : InMux
    port map (
            O => \N__3088\,
            I => \N__3073\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__3083\,
            I => \N__3070\
        );

    \I__658\ : InMux
    port map (
            O => \N__3082\,
            I => \N__3067\
        );

    \I__657\ : InMux
    port map (
            O => \N__3081\,
            I => \N__3062\
        );

    \I__656\ : InMux
    port map (
            O => \N__3080\,
            I => \N__3062\
        );

    \I__655\ : InMux
    port map (
            O => \N__3079\,
            I => \N__3059\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__3076\,
            I => \my_uart.rx_countdown_3_s1_5\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3073\,
            I => \my_uart.rx_countdown_3_s1_5\
        );

    \I__652\ : Odrv12
    port map (
            O => \N__3070\,
            I => \my_uart.rx_countdown_3_s1_5\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__3067\,
            I => \my_uart.rx_countdown_3_s1_5\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__3062\,
            I => \my_uart.rx_countdown_3_s1_5\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__3059\,
            I => \my_uart.rx_countdown_3_s1_5\
        );

    \I__648\ : InMux
    port map (
            O => \N__3046\,
            I => \N__3043\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__3043\,
            I => \my_uart.g0_6_a5_0_3\
        );

    \I__646\ : CascadeMux
    port map (
            O => \N__3040\,
            I => \N__3037\
        );

    \I__645\ : InMux
    port map (
            O => \N__3037\,
            I => \N__3028\
        );

    \I__644\ : InMux
    port map (
            O => \N__3036\,
            I => \N__3028\
        );

    \I__643\ : InMux
    port map (
            O => \N__3035\,
            I => \N__3028\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__3028\,
            I => \my_uart.rx_bits_remainingZ0Z_1\
        );

    \I__641\ : InMux
    port map (
            O => \N__3025\,
            I => \N__3013\
        );

    \I__640\ : InMux
    port map (
            O => \N__3024\,
            I => \N__3013\
        );

    \I__639\ : InMux
    port map (
            O => \N__3023\,
            I => \N__3013\
        );

    \I__638\ : InMux
    port map (
            O => \N__3022\,
            I => \N__3013\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__3013\,
            I => \my_uart.rx_bits_remainingZ0Z_0\
        );

    \I__636\ : InMux
    port map (
            O => \N__3010\,
            I => \N__3007\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__3007\,
            I => \N__3004\
        );

    \I__634\ : Odrv12
    port map (
            O => \N__3004\,
            I => \my_uart.CO1_i\
        );

    \I__633\ : CascadeMux
    port map (
            O => \N__3001\,
            I => \my_uart.CO1_i_cascade_\
        );

    \I__632\ : InMux
    port map (
            O => \N__2998\,
            I => \N__2995\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__2995\,
            I => \N__2990\
        );

    \I__630\ : InMux
    port map (
            O => \N__2994\,
            I => \N__2985\
        );

    \I__629\ : InMux
    port map (
            O => \N__2993\,
            I => \N__2985\
        );

    \I__628\ : Odrv12
    port map (
            O => \N__2990\,
            I => \my_uart.rx_bits_remainingZ0Z_2\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__2985\,
            I => \my_uart.rx_bits_remainingZ0Z_2\
        );

    \I__626\ : CEMux
    port map (
            O => \N__2980\,
            I => \N__2977\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__2977\,
            I => \N__2974\
        );

    \I__624\ : Odrv4
    port map (
            O => \N__2974\,
            I => \my_uart.un1_rx_data_0_sqmuxa_i_i\
        );

    \I__623\ : ClkMux
    port map (
            O => \N__2971\,
            I => \N__2932\
        );

    \I__622\ : ClkMux
    port map (
            O => \N__2970\,
            I => \N__2932\
        );

    \I__621\ : ClkMux
    port map (
            O => \N__2969\,
            I => \N__2932\
        );

    \I__620\ : ClkMux
    port map (
            O => \N__2968\,
            I => \N__2932\
        );

    \I__619\ : ClkMux
    port map (
            O => \N__2967\,
            I => \N__2932\
        );

    \I__618\ : ClkMux
    port map (
            O => \N__2966\,
            I => \N__2932\
        );

    \I__617\ : ClkMux
    port map (
            O => \N__2965\,
            I => \N__2932\
        );

    \I__616\ : ClkMux
    port map (
            O => \N__2964\,
            I => \N__2932\
        );

    \I__615\ : ClkMux
    port map (
            O => \N__2963\,
            I => \N__2932\
        );

    \I__614\ : ClkMux
    port map (
            O => \N__2962\,
            I => \N__2932\
        );

    \I__613\ : ClkMux
    port map (
            O => \N__2961\,
            I => \N__2932\
        );

    \I__612\ : ClkMux
    port map (
            O => \N__2960\,
            I => \N__2932\
        );

    \I__611\ : ClkMux
    port map (
            O => \N__2959\,
            I => \N__2932\
        );

    \I__610\ : GlobalMux
    port map (
            O => \N__2932\,
            I => \N__2929\
        );

    \I__609\ : gio2CtrlBuf
    port map (
            O => \N__2929\,
            I => \CLK_i_c_g\
        );

    \I__608\ : CascadeMux
    port map (
            O => \N__2926\,
            I => \my_uart.m15_e_0_cascade_\
        );

    \I__607\ : CascadeMux
    port map (
            O => \N__2923\,
            I => \my_uart.m15_e_3_cascade_\
        );

    \I__606\ : InMux
    port map (
            O => \N__2920\,
            I => \N__2917\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__2917\,
            I => \my_uart.N_28_mux\
        );

    \I__604\ : InMux
    port map (
            O => \N__2914\,
            I => \N__2911\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__2911\,
            I => \my_uart.N_19_mux_0\
        );

    \I__602\ : InMux
    port map (
            O => \N__2908\,
            I => \N__2905\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__2905\,
            I => \my_uart.m10_e_3\
        );

    \I__600\ : CascadeMux
    port map (
            O => \N__2902\,
            I => \my_uart.N_19_mux_0_cascade_\
        );

    \I__599\ : InMux
    port map (
            O => \N__2899\,
            I => \N__2892\
        );

    \I__598\ : InMux
    port map (
            O => \N__2898\,
            I => \N__2882\
        );

    \I__597\ : CascadeMux
    port map (
            O => \N__2897\,
            I => \N__2878\
        );

    \I__596\ : InMux
    port map (
            O => \N__2896\,
            I => \N__2872\
        );

    \I__595\ : InMux
    port map (
            O => \N__2895\,
            I => \N__2872\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__2892\,
            I => \N__2868\
        );

    \I__593\ : InMux
    port map (
            O => \N__2891\,
            I => \N__2865\
        );

    \I__592\ : CascadeMux
    port map (
            O => \N__2890\,
            I => \N__2859\
        );

    \I__591\ : InMux
    port map (
            O => \N__2889\,
            I => \N__2851\
        );

    \I__590\ : InMux
    port map (
            O => \N__2888\,
            I => \N__2851\
        );

    \I__589\ : InMux
    port map (
            O => \N__2887\,
            I => \N__2851\
        );

    \I__588\ : InMux
    port map (
            O => \N__2886\,
            I => \N__2848\
        );

    \I__587\ : InMux
    port map (
            O => \N__2885\,
            I => \N__2845\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__2882\,
            I => \N__2842\
        );

    \I__585\ : InMux
    port map (
            O => \N__2881\,
            I => \N__2839\
        );

    \I__584\ : InMux
    port map (
            O => \N__2878\,
            I => \N__2834\
        );

    \I__583\ : InMux
    port map (
            O => \N__2877\,
            I => \N__2834\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__2872\,
            I => \N__2831\
        );

    \I__581\ : InMux
    port map (
            O => \N__2871\,
            I => \N__2828\
        );

    \I__580\ : Span4Mux_v
    port map (
            O => \N__2868\,
            I => \N__2823\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__2865\,
            I => \N__2823\
        );

    \I__578\ : InMux
    port map (
            O => \N__2864\,
            I => \N__2818\
        );

    \I__577\ : InMux
    port map (
            O => \N__2863\,
            I => \N__2818\
        );

    \I__576\ : InMux
    port map (
            O => \N__2862\,
            I => \N__2811\
        );

    \I__575\ : InMux
    port map (
            O => \N__2859\,
            I => \N__2811\
        );

    \I__574\ : InMux
    port map (
            O => \N__2858\,
            I => \N__2811\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__2851\,
            I => \my_uart.un1_rx_clk_divider_a\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__2848\,
            I => \my_uart.un1_rx_clk_divider_a\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__2845\,
            I => \my_uart.un1_rx_clk_divider_a\
        );

    \I__570\ : Odrv4
    port map (
            O => \N__2842\,
            I => \my_uart.un1_rx_clk_divider_a\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__2839\,
            I => \my_uart.un1_rx_clk_divider_a\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__2834\,
            I => \my_uart.un1_rx_clk_divider_a\
        );

    \I__567\ : Odrv4
    port map (
            O => \N__2831\,
            I => \my_uart.un1_rx_clk_divider_a\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__2828\,
            I => \my_uart.un1_rx_clk_divider_a\
        );

    \I__565\ : Odrv4
    port map (
            O => \N__2823\,
            I => \my_uart.un1_rx_clk_divider_a\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__2818\,
            I => \my_uart.un1_rx_clk_divider_a\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__2811\,
            I => \my_uart.un1_rx_clk_divider_a\
        );

    \I__562\ : InMux
    port map (
            O => \N__2788\,
            I => \N__2785\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__2785\,
            I => \my_uart.N_27_mux\
        );

    \I__560\ : InMux
    port map (
            O => \N__2782\,
            I => \N__2773\
        );

    \I__559\ : CascadeMux
    port map (
            O => \N__2781\,
            I => \N__2769\
        );

    \I__558\ : InMux
    port map (
            O => \N__2780\,
            I => \N__2763\
        );

    \I__557\ : InMux
    port map (
            O => \N__2779\,
            I => \N__2763\
        );

    \I__556\ : InMux
    port map (
            O => \N__2778\,
            I => \N__2760\
        );

    \I__555\ : InMux
    port map (
            O => \N__2777\,
            I => \N__2757\
        );

    \I__554\ : InMux
    port map (
            O => \N__2776\,
            I => \N__2754\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__2773\,
            I => \N__2751\
        );

    \I__552\ : InMux
    port map (
            O => \N__2772\,
            I => \N__2748\
        );

    \I__551\ : InMux
    port map (
            O => \N__2769\,
            I => \N__2743\
        );

    \I__550\ : InMux
    port map (
            O => \N__2768\,
            I => \N__2743\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__2763\,
            I => \N__2736\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__2760\,
            I => \N__2736\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__2757\,
            I => \N__2736\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__2754\,
            I => \my_uart.rx_countdownZ0Z_5\
        );

    \I__545\ : Odrv4
    port map (
            O => \N__2751\,
            I => \my_uart.rx_countdownZ0Z_5\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__2748\,
            I => \my_uart.rx_countdownZ0Z_5\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__2743\,
            I => \my_uart.rx_countdownZ0Z_5\
        );

    \I__542\ : Odrv4
    port map (
            O => \N__2736\,
            I => \my_uart.rx_countdownZ0Z_5\
        );

    \I__541\ : InMux
    port map (
            O => \N__2725\,
            I => \N__2722\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__2722\,
            I => \my_uart.N_22_mux\
        );

    \I__539\ : CascadeMux
    port map (
            O => \N__2719\,
            I => \my_uart.N_23_mux_cascade_\
        );

    \I__538\ : InMux
    port map (
            O => \N__2716\,
            I => \N__2713\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__2713\,
            I => \my_uart.m7_0_0\
        );

    \I__536\ : InMux
    port map (
            O => \N__2710\,
            I => \N__2707\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__2707\,
            I => \my_uart.g0_6_0_1\
        );

    \I__534\ : CascadeMux
    port map (
            O => \N__2704\,
            I => \my_uart.un1_rx_clk_divider28_i_cascade_\
        );

    \I__533\ : CascadeMux
    port map (
            O => \N__2701\,
            I => \N__2693\
        );

    \I__532\ : CascadeMux
    port map (
            O => \N__2700\,
            I => \N__2690\
        );

    \I__531\ : CascadeMux
    port map (
            O => \N__2699\,
            I => \N__2682\
        );

    \I__530\ : CascadeMux
    port map (
            O => \N__2698\,
            I => \N__2678\
        );

    \I__529\ : SRMux
    port map (
            O => \N__2697\,
            I => \N__2673\
        );

    \I__528\ : InMux
    port map (
            O => \N__2696\,
            I => \N__2662\
        );

    \I__527\ : InMux
    port map (
            O => \N__2693\,
            I => \N__2662\
        );

    \I__526\ : InMux
    port map (
            O => \N__2690\,
            I => \N__2662\
        );

    \I__525\ : InMux
    port map (
            O => \N__2689\,
            I => \N__2662\
        );

    \I__524\ : InMux
    port map (
            O => \N__2688\,
            I => \N__2662\
        );

    \I__523\ : InMux
    port map (
            O => \N__2687\,
            I => \N__2653\
        );

    \I__522\ : InMux
    port map (
            O => \N__2686\,
            I => \N__2653\
        );

    \I__521\ : InMux
    port map (
            O => \N__2685\,
            I => \N__2653\
        );

    \I__520\ : InMux
    port map (
            O => \N__2682\,
            I => \N__2653\
        );

    \I__519\ : InMux
    port map (
            O => \N__2681\,
            I => \N__2650\
        );

    \I__518\ : InMux
    port map (
            O => \N__2678\,
            I => \N__2645\
        );

    \I__517\ : InMux
    port map (
            O => \N__2677\,
            I => \N__2645\
        );

    \I__516\ : CascadeMux
    port map (
            O => \N__2676\,
            I => \N__2642\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__2673\,
            I => \N__2637\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__2662\,
            I => \N__2637\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__2653\,
            I => \N__2634\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__2650\,
            I => \N__2627\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__2645\,
            I => \N__2627\
        );

    \I__510\ : InMux
    port map (
            O => \N__2642\,
            I => \N__2624\
        );

    \I__509\ : Span4Mux_v
    port map (
            O => \N__2637\,
            I => \N__2621\
        );

    \I__508\ : Span4Mux_h
    port map (
            O => \N__2634\,
            I => \N__2618\
        );

    \I__507\ : InMux
    port map (
            O => \N__2633\,
            I => \N__2613\
        );

    \I__506\ : InMux
    port map (
            O => \N__2632\,
            I => \N__2613\
        );

    \I__505\ : Span4Mux_h
    port map (
            O => \N__2627\,
            I => \N__2608\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__2624\,
            I => \N__2608\
        );

    \I__503\ : Odrv4
    port map (
            O => \N__2621\,
            I => \my_uart.rx_clk_divider_0_sqmuxa\
        );

    \I__502\ : Odrv4
    port map (
            O => \N__2618\,
            I => \my_uart.rx_clk_divider_0_sqmuxa\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__2613\,
            I => \my_uart.rx_clk_divider_0_sqmuxa\
        );

    \I__500\ : Odrv4
    port map (
            O => \N__2608\,
            I => \my_uart.rx_clk_divider_0_sqmuxa\
        );

    \I__499\ : InMux
    port map (
            O => \N__2599\,
            I => \N__2596\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__2596\,
            I => \my_uart.m6_0_18_0\
        );

    \I__497\ : CascadeMux
    port map (
            O => \N__2593\,
            I => \N__2589\
        );

    \I__496\ : CascadeMux
    port map (
            O => \N__2592\,
            I => \N__2585\
        );

    \I__495\ : InMux
    port map (
            O => \N__2589\,
            I => \N__2582\
        );

    \I__494\ : InMux
    port map (
            O => \N__2588\,
            I => \N__2577\
        );

    \I__493\ : InMux
    port map (
            O => \N__2585\,
            I => \N__2577\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__2582\,
            I => \N__2574\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__2577\,
            I => \N__2571\
        );

    \I__490\ : Span4Mux_h
    port map (
            O => \N__2574\,
            I => \N__2568\
        );

    \I__489\ : Odrv4
    port map (
            O => \N__2571\,
            I => \my_uart.rx_bits_remainingZ0Z_3\
        );

    \I__488\ : Odrv4
    port map (
            O => \N__2568\,
            I => \my_uart.rx_bits_remainingZ0Z_3\
        );

    \I__487\ : InMux
    port map (
            O => \N__2563\,
            I => \my_uart.rx_countdown_3_cry_3_s1\
        );

    \I__486\ : InMux
    port map (
            O => \N__2560\,
            I => \my_uart.rx_countdown_3_cry_4_s1\
        );

    \I__485\ : CascadeMux
    port map (
            O => \N__2557\,
            I => \N__2554\
        );

    \I__484\ : InMux
    port map (
            O => \N__2554\,
            I => \N__2547\
        );

    \I__483\ : InMux
    port map (
            O => \N__2553\,
            I => \N__2547\
        );

    \I__482\ : InMux
    port map (
            O => \N__2552\,
            I => \N__2544\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__2547\,
            I => \N__2539\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__2544\,
            I => \N__2539\
        );

    \I__479\ : Span4Mux_v
    port map (
            O => \N__2539\,
            I => \N__2534\
        );

    \I__478\ : InMux
    port map (
            O => \N__2538\,
            I => \N__2531\
        );

    \I__477\ : InMux
    port map (
            O => \N__2537\,
            I => \N__2528\
        );

    \I__476\ : Odrv4
    port map (
            O => \N__2534\,
            I => \my_uart.un1_recv_state_8\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__2531\,
            I => \my_uart.un1_recv_state_8\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__2528\,
            I => \my_uart.un1_recv_state_8\
        );

    \I__473\ : InMux
    port map (
            O => \N__2521\,
            I => \N__2518\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__2518\,
            I => \N__2515\
        );

    \I__471\ : Span4Mux_h
    port map (
            O => \N__2515\,
            I => \N__2512\
        );

    \I__470\ : Odrv4
    port map (
            O => \N__2512\,
            I => \my_uart.g0_0_0_a3_3_0\
        );

    \I__469\ : CascadeMux
    port map (
            O => \N__2509\,
            I => \my_uart.N_8_0_cascade_\
        );

    \I__468\ : CascadeMux
    port map (
            O => \N__2506\,
            I => \N__2503\
        );

    \I__467\ : InMux
    port map (
            O => \N__2503\,
            I => \N__2500\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__2500\,
            I => \my_uart.N_18_mux\
        );

    \I__465\ : CascadeMux
    port map (
            O => \N__2497\,
            I => \N__2493\
        );

    \I__464\ : CascadeMux
    port map (
            O => \N__2496\,
            I => \N__2490\
        );

    \I__463\ : InMux
    port map (
            O => \N__2493\,
            I => \N__2485\
        );

    \I__462\ : InMux
    port map (
            O => \N__2490\,
            I => \N__2481\
        );

    \I__461\ : CascadeMux
    port map (
            O => \N__2489\,
            I => \N__2477\
        );

    \I__460\ : CascadeMux
    port map (
            O => \N__2488\,
            I => \N__2474\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__2485\,
            I => \N__2471\
        );

    \I__458\ : CascadeMux
    port map (
            O => \N__2484\,
            I => \N__2466\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__2481\,
            I => \N__2463\
        );

    \I__456\ : InMux
    port map (
            O => \N__2480\,
            I => \N__2458\
        );

    \I__455\ : InMux
    port map (
            O => \N__2477\,
            I => \N__2458\
        );

    \I__454\ : InMux
    port map (
            O => \N__2474\,
            I => \N__2455\
        );

    \I__453\ : Span4Mux_v
    port map (
            O => \N__2471\,
            I => \N__2452\
        );

    \I__452\ : InMux
    port map (
            O => \N__2470\,
            I => \N__2447\
        );

    \I__451\ : InMux
    port map (
            O => \N__2469\,
            I => \N__2447\
        );

    \I__450\ : InMux
    port map (
            O => \N__2466\,
            I => \N__2444\
        );

    \I__449\ : Odrv4
    port map (
            O => \N__2463\,
            I => \my_uart.rx_countdownZ0Z_4\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__2458\,
            I => \my_uart.rx_countdownZ0Z_4\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__2455\,
            I => \my_uart.rx_countdownZ0Z_4\
        );

    \I__446\ : Odrv4
    port map (
            O => \N__2452\,
            I => \my_uart.rx_countdownZ0Z_4\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__2447\,
            I => \my_uart.rx_countdownZ0Z_4\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__2444\,
            I => \my_uart.rx_countdownZ0Z_4\
        );

    \I__443\ : InMux
    port map (
            O => \N__2431\,
            I => \N__2428\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__2428\,
            I => \N__2422\
        );

    \I__441\ : CascadeMux
    port map (
            O => \N__2427\,
            I => \N__2414\
        );

    \I__440\ : InMux
    port map (
            O => \N__2426\,
            I => \N__2409\
        );

    \I__439\ : InMux
    port map (
            O => \N__2425\,
            I => \N__2409\
        );

    \I__438\ : Span4Mux_v
    port map (
            O => \N__2422\,
            I => \N__2406\
        );

    \I__437\ : InMux
    port map (
            O => \N__2421\,
            I => \N__2403\
        );

    \I__436\ : InMux
    port map (
            O => \N__2420\,
            I => \N__2400\
        );

    \I__435\ : InMux
    port map (
            O => \N__2419\,
            I => \N__2397\
        );

    \I__434\ : InMux
    port map (
            O => \N__2418\,
            I => \N__2392\
        );

    \I__433\ : InMux
    port map (
            O => \N__2417\,
            I => \N__2392\
        );

    \I__432\ : InMux
    port map (
            O => \N__2414\,
            I => \N__2389\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__2409\,
            I => \my_uart.rx_countdownZ1Z_1\
        );

    \I__430\ : Odrv4
    port map (
            O => \N__2406\,
            I => \my_uart.rx_countdownZ1Z_1\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__2403\,
            I => \my_uart.rx_countdownZ1Z_1\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__2400\,
            I => \my_uart.rx_countdownZ1Z_1\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__2397\,
            I => \my_uart.rx_countdownZ1Z_1\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__2392\,
            I => \my_uart.rx_countdownZ1Z_1\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__2389\,
            I => \my_uart.rx_countdownZ1Z_1\
        );

    \I__424\ : InMux
    port map (
            O => \N__2374\,
            I => \N__2371\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__2371\,
            I => \N__2363\
        );

    \I__422\ : CascadeMux
    port map (
            O => \N__2370\,
            I => \N__2358\
        );

    \I__421\ : InMux
    port map (
            O => \N__2369\,
            I => \N__2355\
        );

    \I__420\ : InMux
    port map (
            O => \N__2368\,
            I => \N__2352\
        );

    \I__419\ : InMux
    port map (
            O => \N__2367\,
            I => \N__2347\
        );

    \I__418\ : InMux
    port map (
            O => \N__2366\,
            I => \N__2347\
        );

    \I__417\ : Span4Mux_h
    port map (
            O => \N__2363\,
            I => \N__2344\
        );

    \I__416\ : InMux
    port map (
            O => \N__2362\,
            I => \N__2339\
        );

    \I__415\ : InMux
    port map (
            O => \N__2361\,
            I => \N__2339\
        );

    \I__414\ : InMux
    port map (
            O => \N__2358\,
            I => \N__2336\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__2355\,
            I => \my_uart.rx_countdownZ1Z_2\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__2352\,
            I => \my_uart.rx_countdownZ1Z_2\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__2347\,
            I => \my_uart.rx_countdownZ1Z_2\
        );

    \I__410\ : Odrv4
    port map (
            O => \N__2344\,
            I => \my_uart.rx_countdownZ1Z_2\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__2339\,
            I => \my_uart.rx_countdownZ1Z_2\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__2336\,
            I => \my_uart.rx_countdownZ1Z_2\
        );

    \I__407\ : InMux
    port map (
            O => \N__2323\,
            I => \N__2319\
        );

    \I__406\ : InMux
    port map (
            O => \N__2322\,
            I => \N__2315\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__2319\,
            I => \N__2309\
        );

    \I__404\ : InMux
    port map (
            O => \N__2318\,
            I => \N__2306\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__2315\,
            I => \N__2301\
        );

    \I__402\ : InMux
    port map (
            O => \N__2314\,
            I => \N__2298\
        );

    \I__401\ : InMux
    port map (
            O => \N__2313\,
            I => \N__2293\
        );

    \I__400\ : InMux
    port map (
            O => \N__2312\,
            I => \N__2293\
        );

    \I__399\ : Span4Mux_h
    port map (
            O => \N__2309\,
            I => \N__2290\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__2306\,
            I => \N__2287\
        );

    \I__397\ : InMux
    port map (
            O => \N__2305\,
            I => \N__2284\
        );

    \I__396\ : InMux
    port map (
            O => \N__2304\,
            I => \N__2281\
        );

    \I__395\ : Odrv4
    port map (
            O => \N__2301\,
            I => \my_uart.rx_countdownZ1Z_3\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__2298\,
            I => \my_uart.rx_countdownZ1Z_3\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__2293\,
            I => \my_uart.rx_countdownZ1Z_3\
        );

    \I__392\ : Odrv4
    port map (
            O => \N__2290\,
            I => \my_uart.rx_countdownZ1Z_3\
        );

    \I__391\ : Odrv4
    port map (
            O => \N__2287\,
            I => \my_uart.rx_countdownZ1Z_3\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__2284\,
            I => \my_uart.rx_countdownZ1Z_3\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__2281\,
            I => \my_uart.rx_countdownZ1Z_3\
        );

    \I__388\ : CascadeMux
    port map (
            O => \N__2266\,
            I => \my_uart.m10_e_1_cascade_\
        );

    \I__387\ : CascadeMux
    port map (
            O => \N__2263\,
            I => \my_uart.g0_4_a3_3_cascade_\
        );

    \I__386\ : InMux
    port map (
            O => \N__2260\,
            I => \N__2257\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__2257\,
            I => \my_uart.g0_4_a3_4\
        );

    \I__384\ : InMux
    port map (
            O => \N__2254\,
            I => \N__2251\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__2251\,
            I => \my_uart.recv_state_0_sqmuxa_1_0\
        );

    \I__382\ : InMux
    port map (
            O => \N__2248\,
            I => \N__2245\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__2245\,
            I => \my_uart.g0_4_a3_0_2\
        );

    \I__380\ : InMux
    port map (
            O => \N__2242\,
            I => \N__2239\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__2239\,
            I => \my_uart.g0_6_a5_1_0\
        );

    \I__378\ : InMux
    port map (
            O => \N__2236\,
            I => \my_uart.rx_countdown_3_cry_0_s1\
        );

    \I__377\ : InMux
    port map (
            O => \N__2233\,
            I => \my_uart.rx_countdown_3_cry_1_s1\
        );

    \I__376\ : InMux
    port map (
            O => \N__2230\,
            I => \my_uart.rx_countdown_3_cry_2_s1\
        );

    \I__375\ : CascadeMux
    port map (
            O => \N__2227\,
            I => \N__2222\
        );

    \I__374\ : CascadeMux
    port map (
            O => \N__2226\,
            I => \N__2217\
        );

    \I__373\ : InMux
    port map (
            O => \N__2225\,
            I => \N__2210\
        );

    \I__372\ : InMux
    port map (
            O => \N__2222\,
            I => \N__2210\
        );

    \I__371\ : InMux
    port map (
            O => \N__2221\,
            I => \N__2210\
        );

    \I__370\ : InMux
    port map (
            O => \N__2220\,
            I => \N__2204\
        );

    \I__369\ : InMux
    port map (
            O => \N__2217\,
            I => \N__2204\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__2210\,
            I => \N__2194\
        );

    \I__367\ : InMux
    port map (
            O => \N__2209\,
            I => \N__2191\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__2204\,
            I => \N__2188\
        );

    \I__365\ : CascadeMux
    port map (
            O => \N__2203\,
            I => \N__2185\
        );

    \I__364\ : CascadeMux
    port map (
            O => \N__2202\,
            I => \N__2182\
        );

    \I__363\ : CascadeMux
    port map (
            O => \N__2201\,
            I => \N__2179\
        );

    \I__362\ : CascadeMux
    port map (
            O => \N__2200\,
            I => \N__2176\
        );

    \I__361\ : CascadeMux
    port map (
            O => \N__2199\,
            I => \N__2173\
        );

    \I__360\ : CascadeMux
    port map (
            O => \N__2198\,
            I => \N__2170\
        );

    \I__359\ : CascadeMux
    port map (
            O => \N__2197\,
            I => \N__2167\
        );

    \I__358\ : Span4Mux_v
    port map (
            O => \N__2194\,
            I => \N__2164\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__2191\,
            I => \N__2161\
        );

    \I__356\ : Span4Mux_v
    port map (
            O => \N__2188\,
            I => \N__2158\
        );

    \I__355\ : InMux
    port map (
            O => \N__2185\,
            I => \N__2151\
        );

    \I__354\ : InMux
    port map (
            O => \N__2182\,
            I => \N__2151\
        );

    \I__353\ : InMux
    port map (
            O => \N__2179\,
            I => \N__2151\
        );

    \I__352\ : InMux
    port map (
            O => \N__2176\,
            I => \N__2142\
        );

    \I__351\ : InMux
    port map (
            O => \N__2173\,
            I => \N__2142\
        );

    \I__350\ : InMux
    port map (
            O => \N__2170\,
            I => \N__2142\
        );

    \I__349\ : InMux
    port map (
            O => \N__2167\,
            I => \N__2142\
        );

    \I__348\ : Odrv4
    port map (
            O => \N__2164\,
            I => \CONSTANT_ONE_NET\
        );

    \I__347\ : Odrv4
    port map (
            O => \N__2161\,
            I => \CONSTANT_ONE_NET\
        );

    \I__346\ : Odrv4
    port map (
            O => \N__2158\,
            I => \CONSTANT_ONE_NET\
        );

    \I__345\ : LocalMux
    port map (
            O => \N__2151\,
            I => \CONSTANT_ONE_NET\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__2142\,
            I => \CONSTANT_ONE_NET\
        );

    \I__343\ : InMux
    port map (
            O => \N__2131\,
            I => \N__2128\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2128\,
            I => \my_uart.rx_countdown_3_4\
        );

    \I__341\ : CascadeMux
    port map (
            O => \N__2125\,
            I => \my_uart.rx_countdown_3_4_cascade_\
        );

    \I__340\ : InMux
    port map (
            O => \N__2122\,
            I => \N__2119\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__2119\,
            I => \N__2116\
        );

    \I__338\ : Odrv4
    port map (
            O => \N__2116\,
            I => \my_uart.rx_countdown_RNO_4Z0Z_2\
        );

    \I__337\ : InMux
    port map (
            O => \N__2113\,
            I => \N__2110\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2110\,
            I => \my_uart.N_13\
        );

    \I__335\ : InMux
    port map (
            O => \N__2107\,
            I => \N__2101\
        );

    \I__334\ : InMux
    port map (
            O => \N__2106\,
            I => \N__2101\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2101\,
            I => \my_uart.rx_countdown_3_3\
        );

    \I__332\ : InMux
    port map (
            O => \N__2098\,
            I => \N__2095\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__2095\,
            I => \my_uart.G_14_0_a3_0_1\
        );

    \I__330\ : InMux
    port map (
            O => \N__2092\,
            I => \N__2089\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__2089\,
            I => \my_uart.g0_6_0_0\
        );

    \I__328\ : CascadeMux
    port map (
            O => \N__2086\,
            I => \N__2083\
        );

    \I__327\ : InMux
    port map (
            O => \N__2083\,
            I => \N__2080\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__2080\,
            I => \my_uart.g0_4_a3_0_3\
        );

    \I__325\ : CascadeMux
    port map (
            O => \N__2077\,
            I => \my_uart.rx_countdown20_cascade_\
        );

    \I__324\ : InMux
    port map (
            O => \N__2074\,
            I => \N__2071\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__2071\,
            I => \my_uart.un1_recv_state_6\
        );

    \I__322\ : InMux
    port map (
            O => \N__2068\,
            I => \N__2065\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__2065\,
            I => \N__2060\
        );

    \I__320\ : InMux
    port map (
            O => \N__2064\,
            I => \N__2057\
        );

    \I__319\ : CEMux
    port map (
            O => \N__2063\,
            I => \N__2054\
        );

    \I__318\ : Span4Mux_h
    port map (
            O => \N__2060\,
            I => \N__2051\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__2057\,
            I => \my_uart.rx_data_0_sqmuxa\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__2054\,
            I => \my_uart.rx_data_0_sqmuxa\
        );

    \I__315\ : Odrv4
    port map (
            O => \N__2051\,
            I => \my_uart.rx_data_0_sqmuxa\
        );

    \I__314\ : CascadeMux
    port map (
            O => \N__2044\,
            I => \my_uart.N_6_cascade_\
        );

    \I__313\ : InMux
    port map (
            O => \N__2041\,
            I => \N__2038\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__2038\,
            I => \my_uart.un1_rx_clk_divider_a_0\
        );

    \I__311\ : CascadeMux
    port map (
            O => \N__2035\,
            I => \N__2030\
        );

    \I__310\ : InMux
    port map (
            O => \N__2034\,
            I => \N__2027\
        );

    \I__309\ : InMux
    port map (
            O => \N__2033\,
            I => \N__2024\
        );

    \I__308\ : InMux
    port map (
            O => \N__2030\,
            I => \N__2021\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__2027\,
            I => \N__2018\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__2024\,
            I => \my_uart.rx_clk_dividerZ0Z_9\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__2021\,
            I => \my_uart.rx_clk_dividerZ0Z_9\
        );

    \I__304\ : Odrv4
    port map (
            O => \N__2018\,
            I => \my_uart.rx_clk_dividerZ0Z_9\
        );

    \I__303\ : CascadeMux
    port map (
            O => \N__2011\,
            I => \N__2008\
        );

    \I__302\ : InMux
    port map (
            O => \N__2008\,
            I => \N__2005\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__2005\,
            I => \my_uart.un1_rx_clk_divider_a_6\
        );

    \I__300\ : InMux
    port map (
            O => \N__2002\,
            I => \N__1999\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__1999\,
            I => \N__1996\
        );

    \I__298\ : Odrv4
    port map (
            O => \N__1996\,
            I => \my_uart.un1_rx_clk_divider_a_7\
        );

    \I__297\ : CascadeMux
    port map (
            O => \N__1993\,
            I => \my_uart.un1_rx_clk_divider_a_cascade_\
        );

    \I__296\ : InMux
    port map (
            O => \N__1990\,
            I => \N__1987\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__1987\,
            I => \N__1984\
        );

    \I__294\ : Odrv4
    port map (
            O => \N__1984\,
            I => \my_uart.N_5\
        );

    \I__293\ : InMux
    port map (
            O => \N__1981\,
            I => \N__1978\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__1978\,
            I => \my_uart.g0_0_0_a3_0_3\
        );

    \I__291\ : CascadeMux
    port map (
            O => \N__1975\,
            I => \my_uart.g0_6_a5_1_5_cascade_\
        );

    \I__290\ : InMux
    port map (
            O => \N__1972\,
            I => \N__1969\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__1969\,
            I => \my_uart.g0_6_a5_1_4\
        );

    \I__288\ : CascadeMux
    port map (
            O => \N__1966\,
            I => \my_uart.rx_countdown_8_5_cascade_\
        );

    \I__287\ : InMux
    port map (
            O => \N__1963\,
            I => \N__1956\
        );

    \I__286\ : InMux
    port map (
            O => \N__1962\,
            I => \N__1956\
        );

    \I__285\ : InMux
    port map (
            O => \N__1961\,
            I => \N__1953\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__1956\,
            I => \my_uart.rx_clk_dividerZ0Z_8\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__1953\,
            I => \my_uart.rx_clk_dividerZ0Z_8\
        );

    \I__282\ : InMux
    port map (
            O => \N__1948\,
            I => \N__1945\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__1945\,
            I => \my_uart.rx_countdown_RNO_5Z0Z_2\
        );

    \I__280\ : CascadeMux
    port map (
            O => \N__1942\,
            I => \my_uart.rx_countdown_RNO_6Z0Z_2_cascade_\
        );

    \I__279\ : InMux
    port map (
            O => \N__1939\,
            I => \N__1936\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__1936\,
            I => \my_uart.rx_clk_divider_1_cry_6_THRU_CO\
        );

    \I__277\ : InMux
    port map (
            O => \N__1933\,
            I => \N__1928\
        );

    \I__276\ : InMux
    port map (
            O => \N__1932\,
            I => \N__1923\
        );

    \I__275\ : InMux
    port map (
            O => \N__1931\,
            I => \N__1923\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__1928\,
            I => \my_uart.rx_clk_dividerZ0Z_7\
        );

    \I__273\ : LocalMux
    port map (
            O => \N__1923\,
            I => \my_uart.rx_clk_dividerZ0Z_7\
        );

    \I__272\ : InMux
    port map (
            O => \N__1918\,
            I => \N__1915\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__1915\,
            I => \my_uart.rx_clk_divider_1_cry_7_THRU_CO\
        );

    \I__270\ : InMux
    port map (
            O => \N__1912\,
            I => \N__1909\
        );

    \I__269\ : LocalMux
    port map (
            O => \N__1909\,
            I => \my_uart.rx_clk_divider_1_cry_8_THRU_CO\
        );

    \I__268\ : InMux
    port map (
            O => \N__1906\,
            I => \N__1903\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__1903\,
            I => \my_uart.rx_clk_divider_1_cry_1_THRU_CO\
        );

    \I__266\ : InMux
    port map (
            O => \N__1900\,
            I => \N__1895\
        );

    \I__265\ : InMux
    port map (
            O => \N__1899\,
            I => \N__1890\
        );

    \I__264\ : InMux
    port map (
            O => \N__1898\,
            I => \N__1890\
        );

    \I__263\ : LocalMux
    port map (
            O => \N__1895\,
            I => \my_uart.rx_clk_dividerZ0Z_2\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__1890\,
            I => \my_uart.rx_clk_dividerZ0Z_2\
        );

    \I__261\ : InMux
    port map (
            O => \N__1885\,
            I => \N__1882\
        );

    \I__260\ : LocalMux
    port map (
            O => \N__1882\,
            I => \N__1879\
        );

    \I__259\ : Odrv4
    port map (
            O => \N__1879\,
            I => \my_uart.rx_clk_divider_1_cry_2_THRU_CO\
        );

    \I__258\ : InMux
    port map (
            O => \N__1876\,
            I => \N__1873\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__1873\,
            I => \N__1870\
        );

    \I__256\ : Odrv4
    port map (
            O => \N__1870\,
            I => \my_uart.rx_clk_divider_1_cry_3_THRU_CO\
        );

    \I__255\ : InMux
    port map (
            O => \N__1867\,
            I => \N__1864\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__1864\,
            I => \N__1861\
        );

    \I__253\ : Odrv4
    port map (
            O => \N__1861\,
            I => \my_uart.rx_clk_divider_1_cry_5_THRU_CO\
        );

    \I__252\ : InMux
    port map (
            O => \N__1858\,
            I => \N__1855\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__1855\,
            I => \N__1852\
        );

    \I__250\ : Odrv4
    port map (
            O => \N__1852\,
            I => \my_uart.rx_clk_divider_1_cry_4_THRU_CO\
        );

    \I__249\ : InMux
    port map (
            O => \N__1849\,
            I => \N__1845\
        );

    \I__248\ : CascadeMux
    port map (
            O => \N__1848\,
            I => \N__1842\
        );

    \I__247\ : LocalMux
    port map (
            O => \N__1845\,
            I => \N__1838\
        );

    \I__246\ : InMux
    port map (
            O => \N__1842\,
            I => \N__1833\
        );

    \I__245\ : InMux
    port map (
            O => \N__1841\,
            I => \N__1833\
        );

    \I__244\ : Odrv4
    port map (
            O => \N__1838\,
            I => \my_uart.rx_clk_dividerZ0Z_5\
        );

    \I__243\ : LocalMux
    port map (
            O => \N__1833\,
            I => \my_uart.rx_clk_dividerZ0Z_5\
        );

    \I__242\ : CascadeMux
    port map (
            O => \N__1828\,
            I => \N__1824\
        );

    \I__241\ : InMux
    port map (
            O => \N__1827\,
            I => \N__1821\
        );

    \I__240\ : InMux
    port map (
            O => \N__1824\,
            I => \N__1817\
        );

    \I__239\ : LocalMux
    port map (
            O => \N__1821\,
            I => \N__1814\
        );

    \I__238\ : InMux
    port map (
            O => \N__1820\,
            I => \N__1811\
        );

    \I__237\ : LocalMux
    port map (
            O => \N__1817\,
            I => \my_uart.rx_clk_dividerZ0Z_4\
        );

    \I__236\ : Odrv4
    port map (
            O => \N__1814\,
            I => \my_uart.rx_clk_dividerZ0Z_4\
        );

    \I__235\ : LocalMux
    port map (
            O => \N__1811\,
            I => \my_uart.rx_clk_dividerZ0Z_4\
        );

    \I__234\ : InMux
    port map (
            O => \N__1804\,
            I => \N__1800\
        );

    \I__233\ : CascadeMux
    port map (
            O => \N__1803\,
            I => \N__1796\
        );

    \I__232\ : LocalMux
    port map (
            O => \N__1800\,
            I => \N__1793\
        );

    \I__231\ : InMux
    port map (
            O => \N__1799\,
            I => \N__1788\
        );

    \I__230\ : InMux
    port map (
            O => \N__1796\,
            I => \N__1788\
        );

    \I__229\ : Odrv4
    port map (
            O => \N__1793\,
            I => \my_uart.rx_clk_dividerZ0Z_6\
        );

    \I__228\ : LocalMux
    port map (
            O => \N__1788\,
            I => \my_uart.rx_clk_dividerZ0Z_6\
        );

    \I__227\ : InMux
    port map (
            O => \N__1783\,
            I => \N__1780\
        );

    \I__226\ : LocalMux
    port map (
            O => \N__1780\,
            I => \N__1775\
        );

    \I__225\ : InMux
    port map (
            O => \N__1779\,
            I => \N__1770\
        );

    \I__224\ : InMux
    port map (
            O => \N__1778\,
            I => \N__1770\
        );

    \I__223\ : Odrv4
    port map (
            O => \N__1775\,
            I => \my_uart.rx_clk_dividerZ0Z_3\
        );

    \I__222\ : LocalMux
    port map (
            O => \N__1770\,
            I => \my_uart.rx_clk_dividerZ0Z_3\
        );

    \I__221\ : InMux
    port map (
            O => \N__1765\,
            I => \my_uart.rx_clk_divider_1_cry_3\
        );

    \I__220\ : InMux
    port map (
            O => \N__1762\,
            I => \my_uart.rx_clk_divider_1_cry_4\
        );

    \I__219\ : InMux
    port map (
            O => \N__1759\,
            I => \my_uart.rx_clk_divider_1_cry_5\
        );

    \I__218\ : InMux
    port map (
            O => \N__1756\,
            I => \my_uart.rx_clk_divider_1_cry_6\
        );

    \I__217\ : InMux
    port map (
            O => \N__1753\,
            I => \bfn_9_26_0_\
        );

    \I__216\ : InMux
    port map (
            O => \N__1750\,
            I => \my_uart.rx_clk_divider_1_cry_8\
        );

    \I__215\ : InMux
    port map (
            O => \N__1747\,
            I => \my_uart.rx_clk_divider_1_cry_9\
        );

    \I__214\ : InMux
    port map (
            O => \N__1744\,
            I => \N__1740\
        );

    \I__213\ : InMux
    port map (
            O => \N__1743\,
            I => \N__1737\
        );

    \I__212\ : LocalMux
    port map (
            O => \N__1740\,
            I => \my_uart.rx_clk_dividerZ0Z_1\
        );

    \I__211\ : LocalMux
    port map (
            O => \N__1737\,
            I => \my_uart.rx_clk_dividerZ0Z_1\
        );

    \I__210\ : CascadeMux
    port map (
            O => \N__1732\,
            I => \N__1728\
        );

    \I__209\ : InMux
    port map (
            O => \N__1731\,
            I => \N__1725\
        );

    \I__208\ : InMux
    port map (
            O => \N__1728\,
            I => \N__1722\
        );

    \I__207\ : LocalMux
    port map (
            O => \N__1725\,
            I => \my_uart.rx_clk_dividerZ0Z_10\
        );

    \I__206\ : LocalMux
    port map (
            O => \N__1722\,
            I => \my_uart.rx_clk_dividerZ0Z_10\
        );

    \I__205\ : InMux
    port map (
            O => \N__1717\,
            I => \N__1714\
        );

    \I__204\ : LocalMux
    port map (
            O => \N__1714\,
            I => \my_uart.rx_clk_divider_1_cry_0_THRU_CO\
        );

    \I__203\ : InMux
    port map (
            O => \N__1711\,
            I => \N__1706\
        );

    \I__202\ : InMux
    port map (
            O => \N__1710\,
            I => \N__1701\
        );

    \I__201\ : InMux
    port map (
            O => \N__1709\,
            I => \N__1701\
        );

    \I__200\ : LocalMux
    port map (
            O => \N__1706\,
            I => \my_uart.rx_clk_dividerZ1Z_1\
        );

    \I__199\ : LocalMux
    port map (
            O => \N__1701\,
            I => \my_uart.rx_clk_dividerZ1Z_1\
        );

    \I__198\ : IoInMux
    port map (
            O => \N__1696\,
            I => \N__1693\
        );

    \I__197\ : LocalMux
    port map (
            O => \N__1693\,
            I => \N__1690\
        );

    \I__196\ : IoSpan4Mux
    port map (
            O => \N__1690\,
            I => \N__1687\
        );

    \I__195\ : Span4Mux_s1_v
    port map (
            O => \N__1687\,
            I => \N__1684\
        );

    \I__194\ : Span4Mux_v
    port map (
            O => \N__1684\,
            I => \N__1680\
        );

    \I__193\ : InMux
    port map (
            O => \N__1683\,
            I => \N__1677\
        );

    \I__192\ : Odrv4
    port map (
            O => \N__1680\,
            I => \LED_o_c_7\
        );

    \I__191\ : LocalMux
    port map (
            O => \N__1677\,
            I => \LED_o_c_7\
        );

    \I__190\ : IoInMux
    port map (
            O => \N__1672\,
            I => \N__1669\
        );

    \I__189\ : LocalMux
    port map (
            O => \N__1669\,
            I => \N__1666\
        );

    \I__188\ : Span4Mux_s2_v
    port map (
            O => \N__1666\,
            I => \N__1663\
        );

    \I__187\ : Span4Mux_h
    port map (
            O => \N__1663\,
            I => \N__1659\
        );

    \I__186\ : InMux
    port map (
            O => \N__1662\,
            I => \N__1656\
        );

    \I__185\ : Odrv4
    port map (
            O => \N__1659\,
            I => \LED_o_c_6\
        );

    \I__184\ : LocalMux
    port map (
            O => \N__1656\,
            I => \LED_o_c_6\
        );

    \I__183\ : IoInMux
    port map (
            O => \N__1651\,
            I => \N__1648\
        );

    \I__182\ : LocalMux
    port map (
            O => \N__1648\,
            I => \N__1645\
        );

    \I__181\ : IoSpan4Mux
    port map (
            O => \N__1645\,
            I => \N__1642\
        );

    \I__180\ : Span4Mux_s2_v
    port map (
            O => \N__1642\,
            I => \N__1638\
        );

    \I__179\ : InMux
    port map (
            O => \N__1641\,
            I => \N__1635\
        );

    \I__178\ : Odrv4
    port map (
            O => \N__1638\,
            I => \LED_o_c_3\
        );

    \I__177\ : LocalMux
    port map (
            O => \N__1635\,
            I => \LED_o_c_3\
        );

    \I__176\ : IoInMux
    port map (
            O => \N__1630\,
            I => \N__1627\
        );

    \I__175\ : LocalMux
    port map (
            O => \N__1627\,
            I => \N__1624\
        );

    \I__174\ : IoSpan4Mux
    port map (
            O => \N__1624\,
            I => \N__1621\
        );

    \I__173\ : Span4Mux_s2_v
    port map (
            O => \N__1621\,
            I => \N__1617\
        );

    \I__172\ : InMux
    port map (
            O => \N__1620\,
            I => \N__1614\
        );

    \I__171\ : Odrv4
    port map (
            O => \N__1617\,
            I => \LED_o_c_2\
        );

    \I__170\ : LocalMux
    port map (
            O => \N__1614\,
            I => \LED_o_c_2\
        );

    \I__169\ : IoInMux
    port map (
            O => \N__1609\,
            I => \N__1606\
        );

    \I__168\ : LocalMux
    port map (
            O => \N__1606\,
            I => \N__1603\
        );

    \I__167\ : Span4Mux_s1_v
    port map (
            O => \N__1603\,
            I => \N__1600\
        );

    \I__166\ : Span4Mux_v
    port map (
            O => \N__1600\,
            I => \N__1596\
        );

    \I__165\ : InMux
    port map (
            O => \N__1599\,
            I => \N__1593\
        );

    \I__164\ : Odrv4
    port map (
            O => \N__1596\,
            I => \LED_o_c_1\
        );

    \I__163\ : LocalMux
    port map (
            O => \N__1593\,
            I => \LED_o_c_1\
        );

    \I__162\ : IoInMux
    port map (
            O => \N__1588\,
            I => \N__1585\
        );

    \I__161\ : LocalMux
    port map (
            O => \N__1585\,
            I => \N__1582\
        );

    \I__160\ : Span4Mux_s2_v
    port map (
            O => \N__1582\,
            I => \N__1579\
        );

    \I__159\ : Span4Mux_h
    port map (
            O => \N__1579\,
            I => \N__1575\
        );

    \I__158\ : InMux
    port map (
            O => \N__1578\,
            I => \N__1572\
        );

    \I__157\ : Odrv4
    port map (
            O => \N__1575\,
            I => \LED_o_c_5\
        );

    \I__156\ : LocalMux
    port map (
            O => \N__1572\,
            I => \LED_o_c_5\
        );

    \I__155\ : IoInMux
    port map (
            O => \N__1567\,
            I => \N__1564\
        );

    \I__154\ : LocalMux
    port map (
            O => \N__1564\,
            I => \N__1561\
        );

    \I__153\ : Span12Mux_s5_v
    port map (
            O => \N__1561\,
            I => \N__1557\
        );

    \I__152\ : InMux
    port map (
            O => \N__1560\,
            I => \N__1554\
        );

    \I__151\ : Odrv12
    port map (
            O => \N__1557\,
            I => \LED_o_c_4\
        );

    \I__150\ : LocalMux
    port map (
            O => \N__1554\,
            I => \LED_o_c_4\
        );

    \I__149\ : InMux
    port map (
            O => \N__1549\,
            I => \my_uart.rx_clk_divider_1_cry_0\
        );

    \I__148\ : InMux
    port map (
            O => \N__1546\,
            I => \my_uart.rx_clk_divider_1_cry_1\
        );

    \I__147\ : InMux
    port map (
            O => \N__1543\,
            I => \my_uart.rx_clk_divider_1_cry_2\
        );

    \I__146\ : InMux
    port map (
            O => \N__1540\,
            I => \N__1537\
        );

    \I__145\ : LocalMux
    port map (
            O => \N__1537\,
            I => \my_uart.rx_bits_remaining_6_0_3\
        );

    \I__144\ : CascadeMux
    port map (
            O => \N__1534\,
            I => \my_uart.g0_0_0_a3_3_cascade_\
        );

    \I__143\ : CascadeMux
    port map (
            O => \N__1531\,
            I => \my_uart.N_4_cascade_\
        );

    \I__142\ : InMux
    port map (
            O => \N__1528\,
            I => \N__1525\
        );

    \I__141\ : LocalMux
    port map (
            O => \N__1525\,
            I => \N__1522\
        );

    \I__140\ : Odrv4
    port map (
            O => \N__1522\,
            I => \my_uart.g0_0\
        );

    \I__139\ : InMux
    port map (
            O => \N__1519\,
            I => \N__1516\
        );

    \I__138\ : LocalMux
    port map (
            O => \N__1516\,
            I => \my_uart.g0_0_0_a3_4\
        );

    \I__137\ : IoInMux
    port map (
            O => \N__1513\,
            I => \N__1510\
        );

    \I__136\ : LocalMux
    port map (
            O => \N__1510\,
            I => \N__1507\
        );

    \I__135\ : Odrv12
    port map (
            O => \N__1507\,
            I => \LED_o_c_0\
        );

    \I__134\ : CascadeMux
    port map (
            O => \N__1504\,
            I => \my_uart.recv_state_0_sqmuxa_1_cascade_\
        );

    \I__133\ : CascadeMux
    port map (
            O => \N__1501\,
            I => \N__1498\
        );

    \I__132\ : InMux
    port map (
            O => \N__1498\,
            I => \N__1495\
        );

    \I__131\ : LocalMux
    port map (
            O => \N__1495\,
            I => \N__1492\
        );

    \I__130\ : Odrv4
    port map (
            O => \N__1492\,
            I => \my_uart.g0_2\
        );

    \I__129\ : CascadeMux
    port map (
            O => \N__1489\,
            I => \my_uart.g0_0_0_a3_0_0_cascade_\
        );

    \I__128\ : InMux
    port map (
            O => \N__1486\,
            I => \N__1483\
        );

    \I__127\ : LocalMux
    port map (
            O => \N__1483\,
            I => \my_uart.g0_0_0_a3_0_4\
        );

    \IN_MUX_bfv_9_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_25_0_\
        );

    \IN_MUX_bfv_9_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \my_uart.rx_clk_divider_1_cry_7\,
            carryinitout => \bfn_9_26_0_\
        );

    \IN_MUX_bfv_11_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_26_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \my_uart.rx_bits_remaining_RNO_0_3_LC_7_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__1486\,
            in1 => \N__2899\,
            in2 => \N__1501\,
            in3 => \N__1519\,
            lcout => OPEN,
            ltout => \my_uart.recv_state_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_bits_remaining_3_LC_7_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100111010"
        )
    port map (
            in0 => \N__2588\,
            in1 => \N__1540\,
            in2 => \N__1504\,
            in3 => \N__2064\,
            lcout => \my_uart.rx_bits_remainingZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2959\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_bits_remaining_RNO_4_3_LC_7_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__3567\,
            in1 => \N__3305\,
            in2 => \N__3841\,
            in3 => \N__3454\,
            lcout => \my_uart.g0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_bits_remaining_RNO_5_3_LC_7_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2323\,
            in1 => \N__2374\,
            in2 => \N__2497\,
            in3 => \N__3667\,
            lcout => OPEN,
            ltout => \my_uart.g0_0_0_a3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_bits_remaining_RNO_2_3_LC_7_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000010000"
        )
    port map (
            in0 => \N__2431\,
            in1 => \N__2782\,
            in2 => \N__1489\,
            in3 => \_gnd_net_\,
            lcout => \my_uart.g0_0_0_a3_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_bits_remaining_RNO_1_3_LC_7_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000000101"
        )
    port map (
            in0 => \N__3306\,
            in1 => \N__2998\,
            in2 => \N__2592\,
            in3 => \N__3010\,
            lcout => \my_uart.rx_bits_remaining_6_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_RNIH36N1_0_LC_7_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__3190\,
            in1 => \N__3666\,
            in2 => \N__3367\,
            in3 => \N__3718\,
            lcout => OPEN,
            ltout => \my_uart.g0_0_0_a3_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_RNIPOKB5_0_LC_7_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__3091\,
            in1 => \N__3133\,
            in2 => \N__1534\,
            in3 => \N__2891\,
            lcout => OPEN,
            ltout => \my_uart.N_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNI4O0M9_2_LC_7_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000000"
        )
    port map (
            in0 => \N__1990\,
            in1 => \N__3568\,
            in2 => \N__1531\,
            in3 => \N__1528\,
            lcout => \my_uart.rx_data_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNIF559_1_LC_7_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3310\,
            in2 => \_gnd_net_\,
            in3 => \N__3460\,
            lcout => \my_uart.g0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_bits_remaining_RNO_3_3_LC_7_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__3090\,
            in1 => \N__3132\,
            in2 => \_gnd_net_\,
            in3 => \N__2521\,
            lcout => \my_uart.g0_0_0_a3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_data_0_LC_7_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1599\,
            lcout => \LED_o_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2960\,
            ce => \N__2063\,
            sr => \_gnd_net_\
        );

    \my_uart.rx_data_7_LC_7_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__3834\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \LED_o_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2960\,
            ce => \N__2063\,
            sr => \_gnd_net_\
        );

    \my_uart.rx_data_5_LC_7_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1662\,
            lcout => \LED_o_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2960\,
            ce => \N__2063\,
            sr => \_gnd_net_\
        );

    \my_uart.rx_data_2_LC_7_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1641\,
            lcout => \LED_o_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2960\,
            ce => \N__2063\,
            sr => \_gnd_net_\
        );

    \my_uart.rx_data_6_LC_7_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1683\,
            lcout => \LED_o_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2960\,
            ce => \N__2063\,
            sr => \_gnd_net_\
        );

    \my_uart.rx_data_3_LC_7_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1560\,
            lcout => \LED_o_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2960\,
            ce => \N__2063\,
            sr => \_gnd_net_\
        );

    \my_uart.rx_data_1_LC_7_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1620\,
            lcout => \LED_o_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2960\,
            ce => \N__2063\,
            sr => \_gnd_net_\
        );

    \my_uart.rx_data_4_LC_7_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1578\,
            lcout => \LED_o_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2960\,
            ce => \N__2063\,
            sr => \_gnd_net_\
        );

    \my_uart.rx_clk_divider_0_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__2681\,
            in1 => \N__1744\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \my_uart.rx_clk_dividerZ0Z_1\,
            ltout => OPEN,
            carryin => \bfn_9_25_0_\,
            carryout => \my_uart.rx_clk_divider_1_cry_0\,
            clk => \N__2961\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1711\,
            in2 => \N__2197\,
            in3 => \N__1549\,
            lcout => \my_uart.rx_clk_divider_1_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \my_uart.rx_clk_divider_1_cry_0\,
            carryout => \my_uart.rx_clk_divider_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1900\,
            in2 => \N__2201\,
            in3 => \N__1546\,
            lcout => \my_uart.rx_clk_divider_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \my_uart.rx_clk_divider_1_cry_1\,
            carryout => \my_uart.rx_clk_divider_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_clk_divider_1_cry_2_THRU_LUT4_0_LC_9_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1783\,
            in2 => \N__2198\,
            in3 => \N__1543\,
            lcout => \my_uart.rx_clk_divider_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \my_uart.rx_clk_divider_1_cry_2\,
            carryout => \my_uart.rx_clk_divider_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_9_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1827\,
            in2 => \N__2202\,
            in3 => \N__1765\,
            lcout => \my_uart.rx_clk_divider_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \my_uart.rx_clk_divider_1_cry_3\,
            carryout => \my_uart.rx_clk_divider_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_clk_divider_1_cry_4_THRU_LUT4_0_LC_9_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1849\,
            in2 => \N__2199\,
            in3 => \N__1762\,
            lcout => \my_uart.rx_clk_divider_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \my_uart.rx_clk_divider_1_cry_4\,
            carryout => \my_uart.rx_clk_divider_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_clk_divider_1_cry_5_THRU_LUT4_0_LC_9_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1804\,
            in2 => \N__2203\,
            in3 => \N__1759\,
            lcout => \my_uart.rx_clk_divider_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \my_uart.rx_clk_divider_1_cry_5\,
            carryout => \my_uart.rx_clk_divider_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_9_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1933\,
            in2 => \N__2200\,
            in3 => \N__1756\,
            lcout => \my_uart.rx_clk_divider_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \my_uart.rx_clk_divider_1_cry_6\,
            carryout => \my_uart.rx_clk_divider_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_9_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1962\,
            in2 => \N__2226\,
            in3 => \N__1753\,
            lcout => \my_uart.rx_clk_divider_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_9_26_0_\,
            carryout => \my_uart.rx_clk_divider_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_9_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2220\,
            in2 => \N__2035\,
            in3 => \N__1750\,
            lcout => \my_uart.rx_clk_divider_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \my_uart.rx_clk_divider_1_cry_8\,
            carryout => \my_uart.rx_clk_divider_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_clk_divider_10_LC_9_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__1731\,
            in1 => \N__2688\,
            in2 => \_gnd_net_\,
            in3 => \N__1747\,
            lcout => \my_uart.rx_clk_dividerZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2963\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_clk_divider_RNIKT1U_10_LC_9_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__1898\,
            in1 => \N__1743\,
            in2 => \N__1732\,
            in3 => \N__1709\,
            lcout => \my_uart.un1_rx_clk_divider_a_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_clk_divider_1_LC_9_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__1710\,
            in1 => \N__1717\,
            in2 => \_gnd_net_\,
            in3 => \N__2689\,
            lcout => \my_uart.rx_clk_dividerZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2963\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_clk_divider_8_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111001"
        )
    port map (
            in0 => \N__1963\,
            in1 => \N__1918\,
            in2 => \N__2701\,
            in3 => \N__2885\,
            lcout => \my_uart.rx_clk_dividerZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2963\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_clk_divider_9_LC_9_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__2033\,
            in1 => \N__2696\,
            in2 => \_gnd_net_\,
            in3 => \N__1912\,
            lcout => \my_uart.rx_clk_dividerZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2963\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_clk_divider_2_LC_9_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000101"
        )
    port map (
            in0 => \N__1899\,
            in1 => \_gnd_net_\,
            in2 => \N__2700\,
            in3 => \N__1906\,
            lcout => \my_uart.rx_clk_dividerZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2963\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_clk_divider_3_LC_9_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111001"
        )
    port map (
            in0 => \N__1779\,
            in1 => \N__1885\,
            in2 => \N__2699\,
            in3 => \N__2887\,
            lcout => \my_uart.rx_clk_dividerZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2965\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_clk_divider_4_LC_9_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101011"
        )
    port map (
            in0 => \N__2888\,
            in1 => \N__1876\,
            in2 => \N__1828\,
            in3 => \N__2685\,
            lcout => \my_uart.rx_clk_dividerZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2965\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_clk_divider_6_LC_9_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__2687\,
            in1 => \N__1867\,
            in2 => \_gnd_net_\,
            in3 => \N__1799\,
            lcout => \my_uart.rx_clk_dividerZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2965\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_clk_divider_5_LC_9_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011101111"
        )
    port map (
            in0 => \N__2889\,
            in1 => \N__2686\,
            in2 => \N__1848\,
            in3 => \N__1858\,
            lcout => \my_uart.rx_clk_dividerZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2965\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_clk_divider_RNIIMPV_3_LC_9_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__1841\,
            in1 => \N__1820\,
            in2 => \N__1803\,
            in3 => \N__1778\,
            lcout => \my_uart.un1_rx_clk_divider_a_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_RNO_5_2_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2419\,
            in2 => \_gnd_net_\,
            in3 => \N__2768\,
            lcout => \my_uart.rx_countdown_RNO_5Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_RNO_0_5_LC_10_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__3081\,
            in1 => \N__2537\,
            in2 => \N__2781\,
            in3 => \N__2864\,
            lcout => OPEN,
            ltout => \my_uart.rx_countdown_8_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_5_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__2677\,
            in1 => \_gnd_net_\,
            in2 => \N__1966\,
            in3 => \_gnd_net_\,
            lcout => \my_uart.rx_countdownZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2962\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_clk_divider_RNIF1TF_7_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1961\,
            in2 => \_gnd_net_\,
            in3 => \N__1931\,
            lcout => \my_uart.un1_rx_clk_divider_a_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_RNO_6_2_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3080\,
            in2 => \_gnd_net_\,
            in3 => \N__3358\,
            lcout => OPEN,
            ltout => \my_uart.rx_countdown_RNO_6Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_RNO_4_2_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111011101"
        )
    port map (
            in0 => \N__1948\,
            in1 => \N__2863\,
            in2 => \N__1942\,
            in3 => \N__3656\,
            lcout => \my_uart.rx_countdown_RNO_4Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_clk_divider_7_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000101"
        )
    port map (
            in0 => \N__1932\,
            in1 => \_gnd_net_\,
            in2 => \N__2698\,
            in3 => \N__1939\,
            lcout => \my_uart.rx_clk_dividerZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2962\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_RNIDTTP_2_LC_10_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2318\,
            in1 => \N__2369\,
            in2 => \N__2496\,
            in3 => \N__3655\,
            lcout => \my_uart.g0_4_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_1_LC_10_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__2426\,
            in1 => \N__2552\,
            in2 => \N__2897\,
            in3 => \N__3361\,
            lcout => \my_uart.rx_countdownZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2964\,
            ce => 'H',
            sr => \N__2697\
        );

    \my_uart.rx_countdown_RNO_0_2_LC_10_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2367\,
            in1 => \N__2877\,
            in2 => \_gnd_net_\,
            in3 => \N__3188\,
            lcout => OPEN,
            ltout => \my_uart.N_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_2_LC_10_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101000"
        )
    port map (
            in0 => \N__3727\,
            in1 => \N__2068\,
            in2 => \N__2044\,
            in3 => \N__2113\,
            lcout => \my_uart.rx_countdownZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2964\,
            ce => 'H',
            sr => \N__2697\
        );

    \my_uart.rx_clk_divider_RNIU7NL2_9_LC_10_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__2041\,
            in1 => \N__2034\,
            in2 => \N__2011\,
            in3 => \N__2002\,
            lcout => \my_uart.un1_rx_clk_divider_a\,
            ltout => \my_uart.un1_rx_clk_divider_a_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_RNIJ5KS3_5_LC_10_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__2776\,
            in1 => \N__1981\,
            in2 => \N__1993\,
            in3 => \N__2425\,
            lcout => \my_uart.N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_RNIDTTP_0_2_LC_10_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2305\,
            in1 => \N__2366\,
            in2 => \N__2488\,
            in3 => \N__3654\,
            lcout => \my_uart.g0_0_0_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNO_6_0_LC_10_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__3421\,
            in1 => \N__2242\,
            in2 => \N__3304\,
            in3 => \N__2778\,
            lcout => OPEN,
            ltout => \my_uart.g0_6_a5_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNO_1_0_LC_10_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__2862\,
            in1 => \N__1972\,
            in2 => \N__1975\,
            in3 => \N__2092\,
            lcout => \my_uart.g0_6_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_4_LC_10_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__2131\,
            in1 => \_gnd_net_\,
            in2 => \N__2557\,
            in3 => \N__2633\,
            lcout => \my_uart.rx_countdownZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2966\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNO_5_0_LC_10_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2368\,
            in1 => \N__2312\,
            in2 => \N__2489\,
            in3 => \N__2420\,
            lcout => \my_uart.g0_6_a5_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_3_LC_10_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__2553\,
            in1 => \N__2632\,
            in2 => \_gnd_net_\,
            in3 => \N__2107\,
            lcout => \my_uart.rx_countdownZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2966\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_RNINCD63_4_LC_10_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__2480\,
            in1 => \_gnd_net_\,
            in2 => \N__2890\,
            in3 => \N__3130\,
            lcout => \my_uart.rx_countdown_3_4\,
            ltout => \my_uart.rx_countdown_3_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_RNO_2_2_LC_10_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__2098\,
            in1 => \N__2106\,
            in2 => \N__2125\,
            in3 => \N__2122\,
            lcout => \my_uart.N_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_RNIK53C3_3_LC_10_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__2858\,
            in1 => \N__2313\,
            in2 => \_gnd_net_\,
            in3 => \N__3714\,
            lcout => \my_uart.rx_countdown_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_RNO_3_2_LC_10_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__3245\,
            in1 => \N__3420\,
            in2 => \N__3832\,
            in3 => \N__3560\,
            lcout => \my_uart.G_14_0_a3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNO_4_0_LC_10_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000001"
        )
    port map (
            in0 => \N__3244\,
            in1 => \N__3419\,
            in2 => \N__3831\,
            in3 => \N__3559\,
            lcout => \my_uart.g0_6_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_RNIEMHI6_2_LC_11_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__2871\,
            in1 => \N__2248\,
            in2 => \N__2086\,
            in3 => \N__2260\,
            lcout => OPEN,
            ltout => \my_uart.rx_countdown20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNIG81F7_1_LC_11_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__2074\,
            in1 => \_gnd_net_\,
            in2 => \N__2077\,
            in3 => \N__2254\,
            lcout => \my_uart.un1_rx_data_0_sqmuxa_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNIOPND_1_1_LC_11_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__3540\,
            in1 => \_gnd_net_\,
            in2 => \N__3459\,
            in3 => \N__3299\,
            lcout => \my_uart.un1_recv_state_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNIOPND_1_LC_11_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__3297\,
            in1 => \N__3447\,
            in2 => \_gnd_net_\,
            in3 => \N__3538\,
            lcout => \my_uart.un1_recv_state_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_RNIH36N1_0_0_LC_11_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__3189\,
            in1 => \N__3647\,
            in2 => \N__3362\,
            in3 => \N__3710\,
            lcout => OPEN,
            ltout => \my_uart.g0_4_a3_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_RNIRGTL2_0_LC_11_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3124\,
            in2 => \N__2263\,
            in3 => \N__3082\,
            lcout => \my_uart.g0_4_a3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNIAONE_1_LC_11_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__3539\,
            in1 => \N__3806\,
            in2 => \N__3458\,
            in3 => \N__3298\,
            lcout => \my_uart.recv_state_0_sqmuxa_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_RNI80VC_5_LC_11_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2772\,
            in2 => \_gnd_net_\,
            in3 => \N__2421\,
            lcout => \my_uart.g0_4_a3_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNO_8_0_LC_11_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3662\,
            in3 => \N__3516\,
            lcout => \my_uart.g0_6_a5_1_0\,
            ltout => OPEN,
            carryin => \bfn_11_26_0_\,
            carryout => \my_uart.rx_countdown_3_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_3_cry_0_s1_c_RNIE18B_LC_11_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2209\,
            in2 => \N__2427\,
            in3 => \N__2236\,
            lcout => \my_uart.rx_countdown_3_s1_1\,
            ltout => OPEN,
            carryin => \my_uart.rx_countdown_3_cry_0_s1\,
            carryout => \my_uart.rx_countdown_3_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_3_cry_1_s1_c_RNIG7IL_LC_11_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2221\,
            in2 => \N__2370\,
            in3 => \N__2233\,
            lcout => \my_uart.rx_countdown_3_s1_2\,
            ltout => OPEN,
            carryin => \my_uart.rx_countdown_3_cry_1_s1\,
            carryout => \my_uart.rx_countdown_3_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_3_cry_2_s1_c_RNIIDSF_LC_11_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2304\,
            in2 => \N__2227\,
            in3 => \N__2230\,
            lcout => \my_uart.rx_countdown_3_s1_3\,
            ltout => OPEN,
            carryin => \my_uart.rx_countdown_3_cry_2_s1\,
            carryout => \my_uart.rx_countdown_3_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_3_cry_3_s1_c_RNIKJ6A_LC_11_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2225\,
            in2 => \N__2484\,
            in3 => \N__2563\,
            lcout => \my_uart.rx_countdown_3_s1_4\,
            ltout => OPEN,
            carryin => \my_uart.rx_countdown_3_cry_3_s1\,
            carryout => \my_uart.rx_countdown_3_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_3_cry_4_s1_c_RNIMPGK_LC_11_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2777\,
            in2 => \_gnd_net_\,
            in3 => \N__2560\,
            lcout => \my_uart.rx_countdown_3_s1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_0_LC_11_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__3646\,
            in1 => \N__2538\,
            in2 => \N__2676\,
            in3 => \N__2886\,
            lcout => \my_uart.rx_countdownZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2967\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_bits_remaining_RNO_6_3_LC_11_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__3178\,
            in1 => \N__3645\,
            in2 => \N__3363\,
            in3 => \N__3709\,
            lcout => \my_uart.g0_0_0_a3_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNO_0_1_LC_11_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__3586\,
            in1 => \N__2881\,
            in2 => \N__2506\,
            in3 => \N__2716\,
            lcout => OPEN,
            ltout => \my_uart.N_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_1_LC_11_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001110111000000"
        )
    port map (
            in0 => \N__3530\,
            in1 => \N__3282\,
            in2 => \N__2509\,
            in3 => \N__3440\,
            lcout => \N_18_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2969\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNO_4_1_LC_11_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__2470\,
            in1 => \N__2314\,
            in2 => \_gnd_net_\,
            in3 => \N__2361\,
            lcout => \my_uart.N_22_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNO_1_1_LC_11_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2418\,
            in1 => \N__2779\,
            in2 => \N__3556\,
            in3 => \N__3659\,
            lcout => \my_uart.N_18_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNO_4_2_LC_11_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__2469\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2417\,
            lcout => OPEN,
            ltout => \my_uart.m10_e_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNO_2_2_LC_11_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__2362\,
            in1 => \N__2322\,
            in2 => \N__2266\,
            in3 => \N__2780\,
            lcout => \my_uart.m10_e_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNO_5_1_LC_11_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__3122\,
            in1 => \N__3186\,
            in2 => \_gnd_net_\,
            in3 => \N__3715\,
            lcout => OPEN,
            ltout => \my_uart.N_23_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNO_3_1_LC_11_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__3833\,
            in1 => \N__2725\,
            in2 => \N__2719\,
            in3 => \N__3660\,
            lcout => \my_uart.m7_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNO_0_0_LC_11_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__2710\,
            in1 => \N__2898\,
            in2 => \N__3142\,
            in3 => \N__3673\,
            lcout => OPEN,
            ltout => \my_uart.un1_rx_clk_divider28_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_0_LC_11_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000111010"
        )
    port map (
            in0 => \N__3274\,
            in1 => \N__2599\,
            in2 => \N__2704\,
            in3 => \N__3466\,
            lcout => my_uart_recv_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2971\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNIAONE_0_1_LC_11_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3272\,
            in1 => \N__3437\,
            in2 => \N__3829\,
            in3 => \N__3554\,
            lcout => \my_uart.rx_clk_divider_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_cnst_2_0__m6_0_18_0_LC_11_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111000110"
        )
    port map (
            in0 => \N__3273\,
            in1 => \N__3438\,
            in2 => \N__3830\,
            in3 => \N__3555\,
            lcout => \my_uart.m6_0_18_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_cnst_2_0__m6_0_18_a4_1_2_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__2993\,
            in1 => \N__3035\,
            in2 => \N__2593\,
            in3 => \N__3022\,
            lcout => \my_uart.m6_0_18_a4_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_bits_remaining_1_LC_12_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010100101"
        )
    port map (
            in0 => \N__3025\,
            in1 => \_gnd_net_\,
            in2 => \N__3040\,
            in3 => \N__3302\,
            lcout => \my_uart.rx_bits_remainingZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2968\,
            ce => \N__2980\,
            sr => \_gnd_net_\
        );

    \my_uart.rx_bits_remaining_0_LC_12_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__3024\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3301\,
            lcout => \my_uart.rx_bits_remainingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2968\,
            ce => \N__2980\,
            sr => \_gnd_net_\
        );

    \my_uart.rx_bits_remaining_RNINFUH_1_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3036\,
            in2 => \_gnd_net_\,
            in3 => \N__3023\,
            lcout => \my_uart.CO1_i\,
            ltout => \my_uart.CO1_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_bits_remaining_2_LC_12_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2994\,
            in2 => \N__3001\,
            in3 => \N__3303\,
            lcout => \my_uart.rx_bits_remainingZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2968\,
            ce => \N__2980\,
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_2_LC_12_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__2788\,
            in1 => \N__2920\,
            in2 => \_gnd_net_\,
            in3 => \N__3661\,
            lcout => my_uart_recv_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2970\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNO_5_2_LC_12_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3354\,
            in2 => \_gnd_net_\,
            in3 => \N__3185\,
            lcout => OPEN,
            ltout => \my_uart.m15_e_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNO_3_2_LC_12_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__3131\,
            in1 => \N__3089\,
            in2 => \N__2926\,
            in3 => \N__3716\,
            lcout => OPEN,
            ltout => \my_uart.m15_e_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNO_1_2_LC_12_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110011001100"
        )
    port map (
            in0 => \N__3736\,
            in1 => \N__2914\,
            in2 => \N__2923\,
            in3 => \N__2896\,
            lcout => \my_uart.N_28_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNIOPND_0_1_LC_12_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011111111"
        )
    port map (
            in0 => \N__3286\,
            in1 => \N__3423\,
            in2 => \_gnd_net_\,
            in3 => \N__3531\,
            lcout => \my_uart.N_19_mux_0\,
            ltout => \my_uart.N_19_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNO_0_2_LC_12_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001110100"
        )
    port map (
            in0 => \N__3735\,
            in1 => \N__2908\,
            in2 => \N__2902\,
            in3 => \N__2895\,
            lcout => \my_uart.N_27_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RS232_RX_i_ibuf_RNIAONE_LC_12_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__3287\,
            in1 => \N__3422\,
            in2 => \N__3828\,
            in3 => \N__3532\,
            lcout => \N_20_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.rx_countdown_RNO_1_2_LC_12_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__3533\,
            in1 => \N__3288\,
            in2 => \_gnd_net_\,
            in3 => \N__3439\,
            lcout => \my_uart.N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNO_3_0_LC_12_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__3658\,
            in1 => \N__3046\,
            in2 => \N__3558\,
            in3 => \N__3717\,
            lcout => \my_uart.g0_6_a5_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNO_2_1_LC_12_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__3088\,
            in1 => \N__3359\,
            in2 => \N__3557\,
            in3 => \N__3657\,
            lcout => \my_uart.N_19_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_cnst_2_0__m6_0_18_a4_1_LC_12_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__3580\,
            in1 => \N__3271\,
            in2 => \_gnd_net_\,
            in3 => \N__3537\,
            lcout => \my_uart.N_217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNO_2_0_LC_12_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110010"
        )
    port map (
            in0 => \N__3436\,
            in1 => \N__3360\,
            in2 => \N__3300\,
            in3 => \N__3187\,
            lcout => \my_uart.g0_6_a5_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \my_uart.recv_state_RNO_7_0_LC_12_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3123\,
            in2 => \_gnd_net_\,
            in3 => \N__3079\,
            lcout => \my_uart.g0_6_a5_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
