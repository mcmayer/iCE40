// ******************************************************************************

// iCEcube Netlister

// Version:            2016.02.27810

// Build Date:         Jan 28 2016 18:04:03

// File Generated:     Jun 5 2016 21:32:19

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "uart_top" view "INTERFACE"

module uart_top (
    LED_o,
    RS232_TX_o,
    CLK_i,
    RSTn_i,
    RS232_RX_i);

    output [7:0] LED_o;
    input RS232_TX_o;
    input CLK_i;
    input RSTn_i;
    input RS232_RX_i;

    wire N__3943;
    wire N__3942;
    wire N__3941;
    wire N__3932;
    wire N__3931;
    wire N__3930;
    wire N__3923;
    wire N__3922;
    wire N__3921;
    wire N__3914;
    wire N__3913;
    wire N__3912;
    wire N__3905;
    wire N__3904;
    wire N__3903;
    wire N__3896;
    wire N__3895;
    wire N__3894;
    wire N__3887;
    wire N__3886;
    wire N__3885;
    wire N__3878;
    wire N__3877;
    wire N__3876;
    wire N__3869;
    wire N__3868;
    wire N__3867;
    wire N__3860;
    wire N__3859;
    wire N__3858;
    wire N__3841;
    wire N__3838;
    wire N__3835;
    wire N__3834;
    wire N__3833;
    wire N__3832;
    wire N__3831;
    wire N__3830;
    wire N__3829;
    wire N__3828;
    wire N__3825;
    wire N__3822;
    wire N__3819;
    wire N__3816;
    wire N__3813;
    wire N__3810;
    wire N__3807;
    wire N__3806;
    wire N__3803;
    wire N__3798;
    wire N__3795;
    wire N__3790;
    wire N__3785;
    wire N__3782;
    wire N__3779;
    wire N__3776;
    wire N__3773;
    wire N__3768;
    wire N__3765;
    wire N__3762;
    wire N__3755;
    wire N__3752;
    wire N__3747;
    wire N__3744;
    wire N__3741;
    wire N__3736;
    wire N__3735;
    wire N__3730;
    wire N__3727;
    wire N__3724;
    wire N__3721;
    wire N__3718;
    wire N__3717;
    wire N__3716;
    wire N__3715;
    wire N__3714;
    wire N__3711;
    wire N__3710;
    wire N__3709;
    wire N__3706;
    wire N__3703;
    wire N__3700;
    wire N__3697;
    wire N__3694;
    wire N__3691;
    wire N__3688;
    wire N__3673;
    wire N__3670;
    wire N__3667;
    wire N__3666;
    wire N__3663;
    wire N__3662;
    wire N__3661;
    wire N__3660;
    wire N__3659;
    wire N__3658;
    wire N__3657;
    wire N__3656;
    wire N__3655;
    wire N__3654;
    wire N__3651;
    wire N__3648;
    wire N__3647;
    wire N__3646;
    wire N__3645;
    wire N__3642;
    wire N__3639;
    wire N__3634;
    wire N__3629;
    wire N__3624;
    wire N__3621;
    wire N__3618;
    wire N__3615;
    wire N__3612;
    wire N__3605;
    wire N__3586;
    wire N__3583;
    wire N__3580;
    wire N__3577;
    wire N__3574;
    wire N__3571;
    wire N__3568;
    wire N__3567;
    wire N__3564;
    wire N__3561;
    wire N__3560;
    wire N__3559;
    wire N__3558;
    wire N__3557;
    wire N__3556;
    wire N__3555;
    wire N__3554;
    wire N__3549;
    wire N__3544;
    wire N__3541;
    wire N__3540;
    wire N__3539;
    wire N__3538;
    wire N__3537;
    wire N__3534;
    wire N__3533;
    wire N__3532;
    wire N__3531;
    wire N__3530;
    wire N__3527;
    wire N__3522;
    wire N__3517;
    wire N__3516;
    wire N__3513;
    wire N__3506;
    wire N__3501;
    wire N__3494;
    wire N__3489;
    wire N__3484;
    wire N__3481;
    wire N__3466;
    wire N__3463;
    wire N__3460;
    wire N__3459;
    wire N__3458;
    wire N__3455;
    wire N__3454;
    wire N__3451;
    wire N__3448;
    wire N__3447;
    wire N__3444;
    wire N__3441;
    wire N__3440;
    wire N__3439;
    wire N__3438;
    wire N__3437;
    wire N__3436;
    wire N__3429;
    wire N__3424;
    wire N__3423;
    wire N__3422;
    wire N__3421;
    wire N__3420;
    wire N__3419;
    wire N__3416;
    wire N__3413;
    wire N__3408;
    wire N__3405;
    wire N__3402;
    wire N__3399;
    wire N__3394;
    wire N__3391;
    wire N__3386;
    wire N__3367;
    wire N__3364;
    wire N__3363;
    wire N__3362;
    wire N__3361;
    wire N__3360;
    wire N__3359;
    wire N__3358;
    wire N__3355;
    wire N__3354;
    wire N__3351;
    wire N__3348;
    wire N__3345;
    wire N__3340;
    wire N__3337;
    wire N__3334;
    wire N__3331;
    wire N__3328;
    wire N__3325;
    wire N__3310;
    wire N__3307;
    wire N__3306;
    wire N__3305;
    wire N__3304;
    wire N__3303;
    wire N__3302;
    wire N__3301;
    wire N__3300;
    wire N__3299;
    wire N__3298;
    wire N__3297;
    wire N__3294;
    wire N__3289;
    wire N__3288;
    wire N__3287;
    wire N__3286;
    wire N__3283;
    wire N__3282;
    wire N__3275;
    wire N__3274;
    wire N__3273;
    wire N__3272;
    wire N__3271;
    wire N__3268;
    wire N__3261;
    wire N__3256;
    wire N__3249;
    wire N__3246;
    wire N__3245;
    wire N__3244;
    wire N__3241;
    wire N__3238;
    wire N__3231;
    wire N__3226;
    wire N__3223;
    wire N__3220;
    wire N__3217;
    wire N__3214;
    wire N__3209;
    wire N__3190;
    wire N__3189;
    wire N__3188;
    wire N__3187;
    wire N__3186;
    wire N__3185;
    wire N__3182;
    wire N__3179;
    wire N__3178;
    wire N__3175;
    wire N__3172;
    wire N__3169;
    wire N__3166;
    wire N__3163;
    wire N__3160;
    wire N__3157;
    wire N__3142;
    wire N__3139;
    wire N__3136;
    wire N__3133;
    wire N__3132;
    wire N__3131;
    wire N__3130;
    wire N__3125;
    wire N__3124;
    wire N__3123;
    wire N__3122;
    wire N__3119;
    wire N__3116;
    wire N__3113;
    wire N__3110;
    wire N__3107;
    wire N__3104;
    wire N__3091;
    wire N__3090;
    wire N__3089;
    wire N__3088;
    wire N__3083;
    wire N__3082;
    wire N__3081;
    wire N__3080;
    wire N__3079;
    wire N__3076;
    wire N__3073;
    wire N__3070;
    wire N__3067;
    wire N__3062;
    wire N__3059;
    wire N__3046;
    wire N__3043;
    wire N__3040;
    wire N__3037;
    wire N__3036;
    wire N__3035;
    wire N__3028;
    wire N__3025;
    wire N__3024;
    wire N__3023;
    wire N__3022;
    wire N__3013;
    wire N__3010;
    wire N__3007;
    wire N__3004;
    wire N__3001;
    wire N__2998;
    wire N__2995;
    wire N__2994;
    wire N__2993;
    wire N__2990;
    wire N__2985;
    wire N__2980;
    wire N__2977;
    wire N__2974;
    wire N__2971;
    wire N__2970;
    wire N__2969;
    wire N__2968;
    wire N__2967;
    wire N__2966;
    wire N__2965;
    wire N__2964;
    wire N__2963;
    wire N__2962;
    wire N__2961;
    wire N__2960;
    wire N__2959;
    wire N__2932;
    wire N__2929;
    wire N__2926;
    wire N__2923;
    wire N__2920;
    wire N__2917;
    wire N__2914;
    wire N__2911;
    wire N__2908;
    wire N__2905;
    wire N__2902;
    wire N__2899;
    wire N__2898;
    wire N__2897;
    wire N__2896;
    wire N__2895;
    wire N__2892;
    wire N__2891;
    wire N__2890;
    wire N__2889;
    wire N__2888;
    wire N__2887;
    wire N__2886;
    wire N__2885;
    wire N__2882;
    wire N__2881;
    wire N__2878;
    wire N__2877;
    wire N__2872;
    wire N__2871;
    wire N__2868;
    wire N__2865;
    wire N__2864;
    wire N__2863;
    wire N__2862;
    wire N__2859;
    wire N__2858;
    wire N__2851;
    wire N__2848;
    wire N__2845;
    wire N__2842;
    wire N__2839;
    wire N__2834;
    wire N__2831;
    wire N__2828;
    wire N__2823;
    wire N__2818;
    wire N__2811;
    wire N__2788;
    wire N__2785;
    wire N__2782;
    wire N__2781;
    wire N__2780;
    wire N__2779;
    wire N__2778;
    wire N__2777;
    wire N__2776;
    wire N__2773;
    wire N__2772;
    wire N__2769;
    wire N__2768;
    wire N__2763;
    wire N__2760;
    wire N__2757;
    wire N__2754;
    wire N__2751;
    wire N__2748;
    wire N__2743;
    wire N__2736;
    wire N__2725;
    wire N__2722;
    wire N__2719;
    wire N__2716;
    wire N__2713;
    wire N__2710;
    wire N__2707;
    wire N__2704;
    wire N__2701;
    wire N__2700;
    wire N__2699;
    wire N__2698;
    wire N__2697;
    wire N__2696;
    wire N__2693;
    wire N__2690;
    wire N__2689;
    wire N__2688;
    wire N__2687;
    wire N__2686;
    wire N__2685;
    wire N__2682;
    wire N__2681;
    wire N__2678;
    wire N__2677;
    wire N__2676;
    wire N__2673;
    wire N__2662;
    wire N__2653;
    wire N__2650;
    wire N__2645;
    wire N__2642;
    wire N__2637;
    wire N__2634;
    wire N__2633;
    wire N__2632;
    wire N__2627;
    wire N__2624;
    wire N__2621;
    wire N__2618;
    wire N__2613;
    wire N__2608;
    wire N__2599;
    wire N__2596;
    wire N__2593;
    wire N__2592;
    wire N__2589;
    wire N__2588;
    wire N__2585;
    wire N__2582;
    wire N__2577;
    wire N__2574;
    wire N__2571;
    wire N__2568;
    wire N__2563;
    wire N__2560;
    wire N__2557;
    wire N__2554;
    wire N__2553;
    wire N__2552;
    wire N__2547;
    wire N__2544;
    wire N__2539;
    wire N__2538;
    wire N__2537;
    wire N__2534;
    wire N__2531;
    wire N__2528;
    wire N__2521;
    wire N__2518;
    wire N__2515;
    wire N__2512;
    wire N__2509;
    wire N__2506;
    wire N__2503;
    wire N__2500;
    wire N__2497;
    wire N__2496;
    wire N__2493;
    wire N__2490;
    wire N__2489;
    wire N__2488;
    wire N__2485;
    wire N__2484;
    wire N__2481;
    wire N__2480;
    wire N__2477;
    wire N__2474;
    wire N__2471;
    wire N__2470;
    wire N__2469;
    wire N__2466;
    wire N__2463;
    wire N__2458;
    wire N__2455;
    wire N__2452;
    wire N__2447;
    wire N__2444;
    wire N__2431;
    wire N__2428;
    wire N__2427;
    wire N__2426;
    wire N__2425;
    wire N__2422;
    wire N__2421;
    wire N__2420;
    wire N__2419;
    wire N__2418;
    wire N__2417;
    wire N__2414;
    wire N__2409;
    wire N__2406;
    wire N__2403;
    wire N__2400;
    wire N__2397;
    wire N__2392;
    wire N__2389;
    wire N__2374;
    wire N__2371;
    wire N__2370;
    wire N__2369;
    wire N__2368;
    wire N__2367;
    wire N__2366;
    wire N__2363;
    wire N__2362;
    wire N__2361;
    wire N__2358;
    wire N__2355;
    wire N__2352;
    wire N__2347;
    wire N__2344;
    wire N__2339;
    wire N__2336;
    wire N__2323;
    wire N__2322;
    wire N__2319;
    wire N__2318;
    wire N__2315;
    wire N__2314;
    wire N__2313;
    wire N__2312;
    wire N__2309;
    wire N__2306;
    wire N__2305;
    wire N__2304;
    wire N__2301;
    wire N__2298;
    wire N__2293;
    wire N__2290;
    wire N__2287;
    wire N__2284;
    wire N__2281;
    wire N__2266;
    wire N__2263;
    wire N__2260;
    wire N__2257;
    wire N__2254;
    wire N__2251;
    wire N__2248;
    wire N__2245;
    wire N__2242;
    wire N__2239;
    wire N__2236;
    wire N__2233;
    wire N__2230;
    wire N__2227;
    wire N__2226;
    wire N__2225;
    wire N__2222;
    wire N__2221;
    wire N__2220;
    wire N__2217;
    wire N__2210;
    wire N__2209;
    wire N__2204;
    wire N__2203;
    wire N__2202;
    wire N__2201;
    wire N__2200;
    wire N__2199;
    wire N__2198;
    wire N__2197;
    wire N__2194;
    wire N__2191;
    wire N__2188;
    wire N__2185;
    wire N__2182;
    wire N__2179;
    wire N__2176;
    wire N__2173;
    wire N__2170;
    wire N__2167;
    wire N__2164;
    wire N__2161;
    wire N__2158;
    wire N__2151;
    wire N__2142;
    wire N__2131;
    wire N__2128;
    wire N__2125;
    wire N__2122;
    wire N__2119;
    wire N__2116;
    wire N__2113;
    wire N__2110;
    wire N__2107;
    wire N__2106;
    wire N__2101;
    wire N__2098;
    wire N__2095;
    wire N__2092;
    wire N__2089;
    wire N__2086;
    wire N__2083;
    wire N__2080;
    wire N__2077;
    wire N__2074;
    wire N__2071;
    wire N__2068;
    wire N__2065;
    wire N__2064;
    wire N__2063;
    wire N__2060;
    wire N__2057;
    wire N__2054;
    wire N__2051;
    wire N__2044;
    wire N__2041;
    wire N__2038;
    wire N__2035;
    wire N__2034;
    wire N__2033;
    wire N__2030;
    wire N__2027;
    wire N__2024;
    wire N__2021;
    wire N__2018;
    wire N__2011;
    wire N__2008;
    wire N__2005;
    wire N__2002;
    wire N__1999;
    wire N__1996;
    wire N__1993;
    wire N__1990;
    wire N__1987;
    wire N__1984;
    wire N__1981;
    wire N__1978;
    wire N__1975;
    wire N__1972;
    wire N__1969;
    wire N__1966;
    wire N__1963;
    wire N__1962;
    wire N__1961;
    wire N__1956;
    wire N__1953;
    wire N__1948;
    wire N__1945;
    wire N__1942;
    wire N__1939;
    wire N__1936;
    wire N__1933;
    wire N__1932;
    wire N__1931;
    wire N__1928;
    wire N__1923;
    wire N__1918;
    wire N__1915;
    wire N__1912;
    wire N__1909;
    wire N__1906;
    wire N__1903;
    wire N__1900;
    wire N__1899;
    wire N__1898;
    wire N__1895;
    wire N__1890;
    wire N__1885;
    wire N__1882;
    wire N__1879;
    wire N__1876;
    wire N__1873;
    wire N__1870;
    wire N__1867;
    wire N__1864;
    wire N__1861;
    wire N__1858;
    wire N__1855;
    wire N__1852;
    wire N__1849;
    wire N__1848;
    wire N__1845;
    wire N__1842;
    wire N__1841;
    wire N__1838;
    wire N__1833;
    wire N__1828;
    wire N__1827;
    wire N__1824;
    wire N__1821;
    wire N__1820;
    wire N__1817;
    wire N__1814;
    wire N__1811;
    wire N__1804;
    wire N__1803;
    wire N__1800;
    wire N__1799;
    wire N__1796;
    wire N__1793;
    wire N__1788;
    wire N__1783;
    wire N__1780;
    wire N__1779;
    wire N__1778;
    wire N__1775;
    wire N__1770;
    wire N__1765;
    wire N__1762;
    wire N__1759;
    wire N__1756;
    wire N__1753;
    wire N__1750;
    wire N__1747;
    wire N__1744;
    wire N__1743;
    wire N__1740;
    wire N__1737;
    wire N__1732;
    wire N__1731;
    wire N__1728;
    wire N__1725;
    wire N__1722;
    wire N__1717;
    wire N__1714;
    wire N__1711;
    wire N__1710;
    wire N__1709;
    wire N__1706;
    wire N__1701;
    wire N__1696;
    wire N__1693;
    wire N__1690;
    wire N__1687;
    wire N__1684;
    wire N__1683;
    wire N__1680;
    wire N__1677;
    wire N__1672;
    wire N__1669;
    wire N__1666;
    wire N__1663;
    wire N__1662;
    wire N__1659;
    wire N__1656;
    wire N__1651;
    wire N__1648;
    wire N__1645;
    wire N__1642;
    wire N__1641;
    wire N__1638;
    wire N__1635;
    wire N__1630;
    wire N__1627;
    wire N__1624;
    wire N__1621;
    wire N__1620;
    wire N__1617;
    wire N__1614;
    wire N__1609;
    wire N__1606;
    wire N__1603;
    wire N__1600;
    wire N__1599;
    wire N__1596;
    wire N__1593;
    wire N__1588;
    wire N__1585;
    wire N__1582;
    wire N__1579;
    wire N__1578;
    wire N__1575;
    wire N__1572;
    wire N__1567;
    wire N__1564;
    wire N__1561;
    wire N__1560;
    wire N__1557;
    wire N__1554;
    wire N__1549;
    wire N__1546;
    wire N__1543;
    wire N__1540;
    wire N__1537;
    wire N__1534;
    wire N__1531;
    wire N__1528;
    wire N__1525;
    wire N__1522;
    wire N__1519;
    wire N__1516;
    wire N__1513;
    wire N__1510;
    wire N__1507;
    wire N__1504;
    wire N__1501;
    wire N__1498;
    wire N__1495;
    wire N__1492;
    wire N__1489;
    wire N__1486;
    wire N__1483;
    wire GNDG0;
    wire VCCG0;
    wire \my_uart.recv_state_0_sqmuxa_1_cascade_ ;
    wire \my_uart.g0_2 ;
    wire \my_uart.g0_0_0_a3_0_0_cascade_ ;
    wire \my_uart.g0_0_0_a3_0_4 ;
    wire \my_uart.rx_bits_remaining_6_0_3 ;
    wire \my_uart.g0_0_0_a3_3_cascade_ ;
    wire \my_uart.N_4_cascade_ ;
    wire \my_uart.g0_0 ;
    wire \my_uart.g0_0_0_a3_4 ;
    wire LED_o_c_0;
    wire LED_o_c_7;
    wire LED_o_c_6;
    wire LED_o_c_3;
    wire LED_o_c_2;
    wire LED_o_c_1;
    wire LED_o_c_5;
    wire LED_o_c_4;
    wire bfn_9_25_0_;
    wire \my_uart.rx_clk_divider_1_cry_0 ;
    wire \my_uart.rx_clk_divider_1_cry_1 ;
    wire \my_uart.rx_clk_divider_1_cry_2 ;
    wire \my_uart.rx_clk_divider_1_cry_3 ;
    wire \my_uart.rx_clk_divider_1_cry_4 ;
    wire \my_uart.rx_clk_divider_1_cry_5 ;
    wire \my_uart.rx_clk_divider_1_cry_6 ;
    wire \my_uart.rx_clk_divider_1_cry_7 ;
    wire bfn_9_26_0_;
    wire \my_uart.rx_clk_divider_1_cry_8 ;
    wire \my_uart.rx_clk_divider_1_cry_9 ;
    wire \my_uart.rx_clk_dividerZ0Z_1 ;
    wire \my_uart.rx_clk_dividerZ0Z_10 ;
    wire \my_uart.rx_clk_divider_1_cry_0_THRU_CO ;
    wire \my_uart.rx_clk_dividerZ1Z_1 ;
    wire \my_uart.rx_clk_divider_1_cry_7_THRU_CO ;
    wire \my_uart.rx_clk_divider_1_cry_8_THRU_CO ;
    wire \my_uart.rx_clk_divider_1_cry_1_THRU_CO ;
    wire \my_uart.rx_clk_dividerZ0Z_2 ;
    wire \my_uart.rx_clk_divider_1_cry_2_THRU_CO ;
    wire \my_uart.rx_clk_divider_1_cry_3_THRU_CO ;
    wire \my_uart.rx_clk_divider_1_cry_5_THRU_CO ;
    wire \my_uart.rx_clk_divider_1_cry_4_THRU_CO ;
    wire \my_uart.rx_clk_dividerZ0Z_5 ;
    wire \my_uart.rx_clk_dividerZ0Z_4 ;
    wire \my_uart.rx_clk_dividerZ0Z_6 ;
    wire \my_uart.rx_clk_dividerZ0Z_3 ;
    wire \my_uart.rx_countdown_8_5_cascade_ ;
    wire \my_uart.rx_clk_dividerZ0Z_8 ;
    wire \my_uart.rx_countdown_RNO_5Z0Z_2 ;
    wire \my_uart.rx_countdown_RNO_6Z0Z_2_cascade_ ;
    wire \my_uart.rx_clk_divider_1_cry_6_THRU_CO ;
    wire \my_uart.rx_clk_dividerZ0Z_7 ;
    wire \my_uart.rx_data_0_sqmuxa ;
    wire \my_uart.N_6_cascade_ ;
    wire \my_uart.un1_rx_clk_divider_a_0 ;
    wire \my_uart.rx_clk_dividerZ0Z_9 ;
    wire \my_uart.un1_rx_clk_divider_a_6 ;
    wire \my_uart.un1_rx_clk_divider_a_7 ;
    wire \my_uart.un1_rx_clk_divider_a_cascade_ ;
    wire \my_uart.N_5 ;
    wire \my_uart.g0_0_0_a3_0_3 ;
    wire \my_uart.g0_6_a5_1_5_cascade_ ;
    wire \my_uart.g0_6_a5_1_4 ;
    wire \my_uart.rx_countdown_3_4 ;
    wire \my_uart.rx_countdown_3_4_cascade_ ;
    wire \my_uart.rx_countdown_RNO_4Z0Z_2 ;
    wire \my_uart.N_13 ;
    wire \my_uart.rx_countdown_3_3 ;
    wire \my_uart.G_14_0_a3_0_1 ;
    wire \my_uart.g0_6_0_0 ;
    wire \my_uart.g0_4_a3_0_3 ;
    wire \my_uart.rx_countdown20_cascade_ ;
    wire \my_uart.un1_recv_state_6 ;
    wire \my_uart.g0_4_a3_3_cascade_ ;
    wire \my_uart.g0_4_a3_4 ;
    wire \my_uart.recv_state_0_sqmuxa_1_0 ;
    wire \my_uart.g0_4_a3_0_2 ;
    wire \my_uart.g0_6_a5_1_0 ;
    wire bfn_11_26_0_;
    wire \my_uart.rx_countdown_3_cry_0_s1 ;
    wire \my_uart.rx_countdown_3_cry_1_s1 ;
    wire \my_uart.rx_countdown_3_cry_2_s1 ;
    wire CONSTANT_ONE_NET;
    wire \my_uart.rx_countdown_3_cry_3_s1 ;
    wire \my_uart.rx_countdown_3_cry_4_s1 ;
    wire \my_uart.un1_recv_state_8 ;
    wire \my_uart.g0_0_0_a3_3_0 ;
    wire \my_uart.N_8_0_cascade_ ;
    wire \my_uart.N_18_mux ;
    wire \my_uart.rx_countdownZ0Z_4 ;
    wire \my_uart.rx_countdownZ1Z_1 ;
    wire \my_uart.rx_countdownZ1Z_2 ;
    wire \my_uart.rx_countdownZ1Z_3 ;
    wire \my_uart.m10_e_1_cascade_ ;
    wire \my_uart.rx_countdownZ0Z_5 ;
    wire \my_uart.N_22_mux ;
    wire \my_uart.N_23_mux_cascade_ ;
    wire \my_uart.m7_0_0 ;
    wire \my_uart.g0_6_0_1 ;
    wire \my_uart.un1_rx_clk_divider28_i_cascade_ ;
    wire \my_uart.rx_clk_divider_0_sqmuxa ;
    wire \my_uart.m6_0_18_0 ;
    wire \my_uart.rx_bits_remainingZ0Z_3 ;
    wire \my_uart.rx_bits_remainingZ0Z_1 ;
    wire \my_uart.rx_bits_remainingZ0Z_0 ;
    wire \my_uart.CO1_i ;
    wire \my_uart.CO1_i_cascade_ ;
    wire \my_uart.rx_bits_remainingZ0Z_2 ;
    wire \my_uart.un1_rx_data_0_sqmuxa_i_i ;
    wire CLK_i_c_g;
    wire \my_uart.m15_e_0_cascade_ ;
    wire \my_uart.m15_e_3_cascade_ ;
    wire \my_uart.N_28_mux ;
    wire \my_uart.N_19_mux_0 ;
    wire \my_uart.m10_e_3 ;
    wire \my_uart.N_19_mux_0_cascade_ ;
    wire \my_uart.un1_rx_clk_divider_a ;
    wire \my_uart.N_27_mux ;
    wire RS232_RX_i_c;
    wire N_20_mux;
    wire \my_uart.N_11 ;
    wire \my_uart.rx_countdown_3_s1_3 ;
    wire \my_uart.g0_6_a5_0_5 ;
    wire \my_uart.rx_countdownZ0Z_3 ;
    wire \my_uart.N_19_mux ;
    wire \my_uart.m6_0_18_a4_1_2 ;
    wire my_uart_recv_state_2;
    wire \my_uart.N_217 ;
    wire N_18_i;
    wire \my_uart.rx_countdown_3_s1_1 ;
    wire my_uart_recv_state_0;
    wire \my_uart.rx_countdown_3_s1_2 ;
    wire \my_uart.g0_6_a5_0_4 ;
    wire \my_uart.rx_countdown_3_s1_4 ;
    wire \my_uart.rx_countdown_3_s1_5 ;
    wire \my_uart.g0_6_a5_0_3 ;
    wire _gnd_net_;

    PRE_IO_GBUF CLK_i_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__3941),
            .GLOBALBUFFEROUTPUT(CLK_i_c_g));
    IO_PAD CLK_i_ibuf_gb_io_iopad (
            .OE(N__3943),
            .DIN(N__3942),
            .DOUT(N__3941),
            .PACKAGEPIN(CLK_i));
    defparam CLK_i_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK_i_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_i_ibuf_gb_io_preio (
            .PADOEN(N__3943),
            .PADOUT(N__3942),
            .PADIN(N__3941),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED_o_obuf_0_iopad (
            .OE(N__3932),
            .DIN(N__3931),
            .DOUT(N__3930),
            .PACKAGEPIN(LED_o[0]));
    defparam LED_o_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam LED_o_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_o_obuf_0_preio (
            .PADOEN(N__3932),
            .PADOUT(N__3931),
            .PADIN(N__3930),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1513),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED_o_obuf_5_iopad (
            .OE(N__3923),
            .DIN(N__3922),
            .DOUT(N__3921),
            .PACKAGEPIN(LED_o[5]));
    defparam LED_o_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam LED_o_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_o_obuf_5_preio (
            .PADOEN(N__3923),
            .PADOUT(N__3922),
            .PADIN(N__3921),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1588),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED_o_obuf_1_iopad (
            .OE(N__3914),
            .DIN(N__3913),
            .DOUT(N__3912),
            .PACKAGEPIN(LED_o[1]));
    defparam LED_o_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam LED_o_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_o_obuf_1_preio (
            .PADOEN(N__3914),
            .PADOUT(N__3913),
            .PADIN(N__3912),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1609),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED_o_obuf_6_iopad (
            .OE(N__3905),
            .DIN(N__3904),
            .DOUT(N__3903),
            .PACKAGEPIN(LED_o[6]));
    defparam LED_o_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam LED_o_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_o_obuf_6_preio (
            .PADOEN(N__3905),
            .PADOUT(N__3904),
            .PADIN(N__3903),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1672),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED_o_obuf_2_iopad (
            .OE(N__3896),
            .DIN(N__3895),
            .DOUT(N__3894),
            .PACKAGEPIN(LED_o[2]));
    defparam LED_o_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam LED_o_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_o_obuf_2_preio (
            .PADOEN(N__3896),
            .PADOUT(N__3895),
            .PADIN(N__3894),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1630),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RS232_RX_i_ibuf_iopad (
            .OE(N__3887),
            .DIN(N__3886),
            .DOUT(N__3885),
            .PACKAGEPIN(RS232_RX_i));
    defparam RS232_RX_i_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RS232_RX_i_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RS232_RX_i_ibuf_preio (
            .PADOEN(N__3887),
            .PADOUT(N__3886),
            .PADIN(N__3885),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RS232_RX_i_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED_o_obuf_7_iopad (
            .OE(N__3878),
            .DIN(N__3877),
            .DOUT(N__3876),
            .PACKAGEPIN(LED_o[7]));
    defparam LED_o_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam LED_o_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_o_obuf_7_preio (
            .PADOEN(N__3878),
            .PADOUT(N__3877),
            .PADIN(N__3876),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1696),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED_o_obuf_3_iopad (
            .OE(N__3869),
            .DIN(N__3868),
            .DOUT(N__3867),
            .PACKAGEPIN(LED_o[3]));
    defparam LED_o_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam LED_o_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_o_obuf_3_preio (
            .PADOEN(N__3869),
            .PADOUT(N__3868),
            .PADIN(N__3867),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1651),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED_o_obuf_4_iopad (
            .OE(N__3860),
            .DIN(N__3859),
            .DOUT(N__3858),
            .PACKAGEPIN(LED_o[4]));
    defparam LED_o_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam LED_o_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_o_obuf_4_preio (
            .PADOEN(N__3860),
            .PADOUT(N__3859),
            .PADIN(N__3858),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1567),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__913 (
            .O(N__3841),
            .I(N__3838));
    InMux I__912 (
            .O(N__3838),
            .I(N__3835));
    LocalMux I__911 (
            .O(N__3835),
            .I(N__3825));
    InMux I__910 (
            .O(N__3834),
            .I(N__3822));
    InMux I__909 (
            .O(N__3833),
            .I(N__3819));
    CascadeMux I__908 (
            .O(N__3832),
            .I(N__3816));
    CascadeMux I__907 (
            .O(N__3831),
            .I(N__3813));
    CascadeMux I__906 (
            .O(N__3830),
            .I(N__3810));
    CascadeMux I__905 (
            .O(N__3829),
            .I(N__3807));
    CascadeMux I__904 (
            .O(N__3828),
            .I(N__3803));
    Span4Mux_v I__903 (
            .O(N__3825),
            .I(N__3798));
    LocalMux I__902 (
            .O(N__3822),
            .I(N__3798));
    LocalMux I__901 (
            .O(N__3819),
            .I(N__3795));
    InMux I__900 (
            .O(N__3816),
            .I(N__3790));
    InMux I__899 (
            .O(N__3813),
            .I(N__3790));
    InMux I__898 (
            .O(N__3810),
            .I(N__3785));
    InMux I__897 (
            .O(N__3807),
            .I(N__3785));
    InMux I__896 (
            .O(N__3806),
            .I(N__3782));
    InMux I__895 (
            .O(N__3803),
            .I(N__3779));
    Span4Mux_v I__894 (
            .O(N__3798),
            .I(N__3776));
    Span4Mux_v I__893 (
            .O(N__3795),
            .I(N__3773));
    LocalMux I__892 (
            .O(N__3790),
            .I(N__3768));
    LocalMux I__891 (
            .O(N__3785),
            .I(N__3768));
    LocalMux I__890 (
            .O(N__3782),
            .I(N__3765));
    LocalMux I__889 (
            .O(N__3779),
            .I(N__3762));
    Span4Mux_h I__888 (
            .O(N__3776),
            .I(N__3755));
    Span4Mux_s3_v I__887 (
            .O(N__3773),
            .I(N__3755));
    Span4Mux_v I__886 (
            .O(N__3768),
            .I(N__3755));
    Sp12to4 I__885 (
            .O(N__3765),
            .I(N__3752));
    Span12Mux_v I__884 (
            .O(N__3762),
            .I(N__3747));
    Sp12to4 I__883 (
            .O(N__3755),
            .I(N__3747));
    Span12Mux_h I__882 (
            .O(N__3752),
            .I(N__3744));
    Span12Mux_h I__881 (
            .O(N__3747),
            .I(N__3741));
    Odrv12 I__880 (
            .O(N__3744),
            .I(RS232_RX_i_c));
    Odrv12 I__879 (
            .O(N__3741),
            .I(RS232_RX_i_c));
    InMux I__878 (
            .O(N__3736),
            .I(N__3730));
    InMux I__877 (
            .O(N__3735),
            .I(N__3730));
    LocalMux I__876 (
            .O(N__3730),
            .I(N_20_mux));
    InMux I__875 (
            .O(N__3727),
            .I(N__3724));
    LocalMux I__874 (
            .O(N__3724),
            .I(N__3721));
    Odrv4 I__873 (
            .O(N__3721),
            .I(\my_uart.N_11 ));
    InMux I__872 (
            .O(N__3718),
            .I(N__3711));
    InMux I__871 (
            .O(N__3717),
            .I(N__3706));
    InMux I__870 (
            .O(N__3716),
            .I(N__3703));
    InMux I__869 (
            .O(N__3715),
            .I(N__3700));
    InMux I__868 (
            .O(N__3714),
            .I(N__3697));
    LocalMux I__867 (
            .O(N__3711),
            .I(N__3694));
    InMux I__866 (
            .O(N__3710),
            .I(N__3691));
    InMux I__865 (
            .O(N__3709),
            .I(N__3688));
    LocalMux I__864 (
            .O(N__3706),
            .I(\my_uart.rx_countdown_3_s1_3 ));
    LocalMux I__863 (
            .O(N__3703),
            .I(\my_uart.rx_countdown_3_s1_3 ));
    LocalMux I__862 (
            .O(N__3700),
            .I(\my_uart.rx_countdown_3_s1_3 ));
    LocalMux I__861 (
            .O(N__3697),
            .I(\my_uart.rx_countdown_3_s1_3 ));
    Odrv12 I__860 (
            .O(N__3694),
            .I(\my_uart.rx_countdown_3_s1_3 ));
    LocalMux I__859 (
            .O(N__3691),
            .I(\my_uart.rx_countdown_3_s1_3 ));
    LocalMux I__858 (
            .O(N__3688),
            .I(\my_uart.rx_countdown_3_s1_3 ));
    InMux I__857 (
            .O(N__3673),
            .I(N__3670));
    LocalMux I__856 (
            .O(N__3670),
            .I(\my_uart.g0_6_a5_0_5 ));
    InMux I__855 (
            .O(N__3667),
            .I(N__3663));
    InMux I__854 (
            .O(N__3666),
            .I(N__3651));
    LocalMux I__853 (
            .O(N__3663),
            .I(N__3648));
    CascadeMux I__852 (
            .O(N__3662),
            .I(N__3642));
    InMux I__851 (
            .O(N__3661),
            .I(N__3639));
    InMux I__850 (
            .O(N__3660),
            .I(N__3634));
    InMux I__849 (
            .O(N__3659),
            .I(N__3634));
    InMux I__848 (
            .O(N__3658),
            .I(N__3629));
    InMux I__847 (
            .O(N__3657),
            .I(N__3629));
    InMux I__846 (
            .O(N__3656),
            .I(N__3624));
    InMux I__845 (
            .O(N__3655),
            .I(N__3624));
    InMux I__844 (
            .O(N__3654),
            .I(N__3621));
    LocalMux I__843 (
            .O(N__3651),
            .I(N__3618));
    Span4Mux_h I__842 (
            .O(N__3648),
            .I(N__3615));
    InMux I__841 (
            .O(N__3647),
            .I(N__3612));
    InMux I__840 (
            .O(N__3646),
            .I(N__3605));
    InMux I__839 (
            .O(N__3645),
            .I(N__3605));
    InMux I__838 (
            .O(N__3642),
            .I(N__3605));
    LocalMux I__837 (
            .O(N__3639),
            .I(\my_uart.rx_countdownZ0Z_3 ));
    LocalMux I__836 (
            .O(N__3634),
            .I(\my_uart.rx_countdownZ0Z_3 ));
    LocalMux I__835 (
            .O(N__3629),
            .I(\my_uart.rx_countdownZ0Z_3 ));
    LocalMux I__834 (
            .O(N__3624),
            .I(\my_uart.rx_countdownZ0Z_3 ));
    LocalMux I__833 (
            .O(N__3621),
            .I(\my_uart.rx_countdownZ0Z_3 ));
    Odrv12 I__832 (
            .O(N__3618),
            .I(\my_uart.rx_countdownZ0Z_3 ));
    Odrv4 I__831 (
            .O(N__3615),
            .I(\my_uart.rx_countdownZ0Z_3 ));
    LocalMux I__830 (
            .O(N__3612),
            .I(\my_uart.rx_countdownZ0Z_3 ));
    LocalMux I__829 (
            .O(N__3605),
            .I(\my_uart.rx_countdownZ0Z_3 ));
    InMux I__828 (
            .O(N__3586),
            .I(N__3583));
    LocalMux I__827 (
            .O(N__3583),
            .I(\my_uart.N_19_mux ));
    InMux I__826 (
            .O(N__3580),
            .I(N__3577));
    LocalMux I__825 (
            .O(N__3577),
            .I(N__3574));
    Span4Mux_h I__824 (
            .O(N__3574),
            .I(N__3571));
    Odrv4 I__823 (
            .O(N__3571),
            .I(\my_uart.m6_0_18_a4_1_2 ));
    InMux I__822 (
            .O(N__3568),
            .I(N__3564));
    InMux I__821 (
            .O(N__3567),
            .I(N__3561));
    LocalMux I__820 (
            .O(N__3564),
            .I(N__3549));
    LocalMux I__819 (
            .O(N__3561),
            .I(N__3549));
    InMux I__818 (
            .O(N__3560),
            .I(N__3544));
    InMux I__817 (
            .O(N__3559),
            .I(N__3544));
    CascadeMux I__816 (
            .O(N__3558),
            .I(N__3541));
    CascadeMux I__815 (
            .O(N__3557),
            .I(N__3534));
    CascadeMux I__814 (
            .O(N__3556),
            .I(N__3527));
    InMux I__813 (
            .O(N__3555),
            .I(N__3522));
    InMux I__812 (
            .O(N__3554),
            .I(N__3522));
    Span4Mux_v I__811 (
            .O(N__3549),
            .I(N__3517));
    LocalMux I__810 (
            .O(N__3544),
            .I(N__3517));
    InMux I__809 (
            .O(N__3541),
            .I(N__3513));
    InMux I__808 (
            .O(N__3540),
            .I(N__3506));
    InMux I__807 (
            .O(N__3539),
            .I(N__3506));
    InMux I__806 (
            .O(N__3538),
            .I(N__3506));
    InMux I__805 (
            .O(N__3537),
            .I(N__3501));
    InMux I__804 (
            .O(N__3534),
            .I(N__3501));
    InMux I__803 (
            .O(N__3533),
            .I(N__3494));
    InMux I__802 (
            .O(N__3532),
            .I(N__3494));
    InMux I__801 (
            .O(N__3531),
            .I(N__3494));
    InMux I__800 (
            .O(N__3530),
            .I(N__3489));
    InMux I__799 (
            .O(N__3527),
            .I(N__3489));
    LocalMux I__798 (
            .O(N__3522),
            .I(N__3484));
    Span4Mux_h I__797 (
            .O(N__3517),
            .I(N__3484));
    InMux I__796 (
            .O(N__3516),
            .I(N__3481));
    LocalMux I__795 (
            .O(N__3513),
            .I(my_uart_recv_state_2));
    LocalMux I__794 (
            .O(N__3506),
            .I(my_uart_recv_state_2));
    LocalMux I__793 (
            .O(N__3501),
            .I(my_uart_recv_state_2));
    LocalMux I__792 (
            .O(N__3494),
            .I(my_uart_recv_state_2));
    LocalMux I__791 (
            .O(N__3489),
            .I(my_uart_recv_state_2));
    Odrv4 I__790 (
            .O(N__3484),
            .I(my_uart_recv_state_2));
    LocalMux I__789 (
            .O(N__3481),
            .I(my_uart_recv_state_2));
    InMux I__788 (
            .O(N__3466),
            .I(N__3463));
    LocalMux I__787 (
            .O(N__3463),
            .I(\my_uart.N_217 ));
    InMux I__786 (
            .O(N__3460),
            .I(N__3455));
    CascadeMux I__785 (
            .O(N__3459),
            .I(N__3451));
    CascadeMux I__784 (
            .O(N__3458),
            .I(N__3448));
    LocalMux I__783 (
            .O(N__3455),
            .I(N__3444));
    InMux I__782 (
            .O(N__3454),
            .I(N__3441));
    InMux I__781 (
            .O(N__3451),
            .I(N__3429));
    InMux I__780 (
            .O(N__3448),
            .I(N__3429));
    InMux I__779 (
            .O(N__3447),
            .I(N__3429));
    Span4Mux_v I__778 (
            .O(N__3444),
            .I(N__3424));
    LocalMux I__777 (
            .O(N__3441),
            .I(N__3424));
    InMux I__776 (
            .O(N__3440),
            .I(N__3416));
    InMux I__775 (
            .O(N__3439),
            .I(N__3413));
    InMux I__774 (
            .O(N__3438),
            .I(N__3408));
    InMux I__773 (
            .O(N__3437),
            .I(N__3408));
    InMux I__772 (
            .O(N__3436),
            .I(N__3405));
    LocalMux I__771 (
            .O(N__3429),
            .I(N__3402));
    Span4Mux_h I__770 (
            .O(N__3424),
            .I(N__3399));
    InMux I__769 (
            .O(N__3423),
            .I(N__3394));
    InMux I__768 (
            .O(N__3422),
            .I(N__3394));
    InMux I__767 (
            .O(N__3421),
            .I(N__3391));
    InMux I__766 (
            .O(N__3420),
            .I(N__3386));
    InMux I__765 (
            .O(N__3419),
            .I(N__3386));
    LocalMux I__764 (
            .O(N__3416),
            .I(N_18_i));
    LocalMux I__763 (
            .O(N__3413),
            .I(N_18_i));
    LocalMux I__762 (
            .O(N__3408),
            .I(N_18_i));
    LocalMux I__761 (
            .O(N__3405),
            .I(N_18_i));
    Odrv4 I__760 (
            .O(N__3402),
            .I(N_18_i));
    Odrv4 I__759 (
            .O(N__3399),
            .I(N_18_i));
    LocalMux I__758 (
            .O(N__3394),
            .I(N_18_i));
    LocalMux I__757 (
            .O(N__3391),
            .I(N_18_i));
    LocalMux I__756 (
            .O(N__3386),
            .I(N_18_i));
    CascadeMux I__755 (
            .O(N__3367),
            .I(N__3364));
    InMux I__754 (
            .O(N__3364),
            .I(N__3355));
    CascadeMux I__753 (
            .O(N__3363),
            .I(N__3351));
    CascadeMux I__752 (
            .O(N__3362),
            .I(N__3348));
    InMux I__751 (
            .O(N__3361),
            .I(N__3345));
    InMux I__750 (
            .O(N__3360),
            .I(N__3340));
    InMux I__749 (
            .O(N__3359),
            .I(N__3340));
    InMux I__748 (
            .O(N__3358),
            .I(N__3337));
    LocalMux I__747 (
            .O(N__3355),
            .I(N__3334));
    InMux I__746 (
            .O(N__3354),
            .I(N__3331));
    InMux I__745 (
            .O(N__3351),
            .I(N__3328));
    InMux I__744 (
            .O(N__3348),
            .I(N__3325));
    LocalMux I__743 (
            .O(N__3345),
            .I(\my_uart.rx_countdown_3_s1_1 ));
    LocalMux I__742 (
            .O(N__3340),
            .I(\my_uart.rx_countdown_3_s1_1 ));
    LocalMux I__741 (
            .O(N__3337),
            .I(\my_uart.rx_countdown_3_s1_1 ));
    Odrv12 I__740 (
            .O(N__3334),
            .I(\my_uart.rx_countdown_3_s1_1 ));
    LocalMux I__739 (
            .O(N__3331),
            .I(\my_uart.rx_countdown_3_s1_1 ));
    LocalMux I__738 (
            .O(N__3328),
            .I(\my_uart.rx_countdown_3_s1_1 ));
    LocalMux I__737 (
            .O(N__3325),
            .I(\my_uart.rx_countdown_3_s1_1 ));
    InMux I__736 (
            .O(N__3310),
            .I(N__3307));
    LocalMux I__735 (
            .O(N__3307),
            .I(N__3294));
    InMux I__734 (
            .O(N__3306),
            .I(N__3289));
    InMux I__733 (
            .O(N__3305),
            .I(N__3289));
    CascadeMux I__732 (
            .O(N__3304),
            .I(N__3283));
    InMux I__731 (
            .O(N__3303),
            .I(N__3275));
    InMux I__730 (
            .O(N__3302),
            .I(N__3275));
    InMux I__729 (
            .O(N__3301),
            .I(N__3275));
    CascadeMux I__728 (
            .O(N__3300),
            .I(N__3268));
    InMux I__727 (
            .O(N__3299),
            .I(N__3261));
    InMux I__726 (
            .O(N__3298),
            .I(N__3261));
    InMux I__725 (
            .O(N__3297),
            .I(N__3261));
    Span4Mux_v I__724 (
            .O(N__3294),
            .I(N__3256));
    LocalMux I__723 (
            .O(N__3289),
            .I(N__3256));
    InMux I__722 (
            .O(N__3288),
            .I(N__3249));
    InMux I__721 (
            .O(N__3287),
            .I(N__3249));
    InMux I__720 (
            .O(N__3286),
            .I(N__3249));
    InMux I__719 (
            .O(N__3283),
            .I(N__3246));
    InMux I__718 (
            .O(N__3282),
            .I(N__3241));
    LocalMux I__717 (
            .O(N__3275),
            .I(N__3238));
    InMux I__716 (
            .O(N__3274),
            .I(N__3231));
    InMux I__715 (
            .O(N__3273),
            .I(N__3231));
    InMux I__714 (
            .O(N__3272),
            .I(N__3231));
    InMux I__713 (
            .O(N__3271),
            .I(N__3226));
    InMux I__712 (
            .O(N__3268),
            .I(N__3226));
    LocalMux I__711 (
            .O(N__3261),
            .I(N__3223));
    Span4Mux_h I__710 (
            .O(N__3256),
            .I(N__3220));
    LocalMux I__709 (
            .O(N__3249),
            .I(N__3217));
    LocalMux I__708 (
            .O(N__3246),
            .I(N__3214));
    InMux I__707 (
            .O(N__3245),
            .I(N__3209));
    InMux I__706 (
            .O(N__3244),
            .I(N__3209));
    LocalMux I__705 (
            .O(N__3241),
            .I(my_uart_recv_state_0));
    Odrv4 I__704 (
            .O(N__3238),
            .I(my_uart_recv_state_0));
    LocalMux I__703 (
            .O(N__3231),
            .I(my_uart_recv_state_0));
    LocalMux I__702 (
            .O(N__3226),
            .I(my_uart_recv_state_0));
    Odrv4 I__701 (
            .O(N__3223),
            .I(my_uart_recv_state_0));
    Odrv4 I__700 (
            .O(N__3220),
            .I(my_uart_recv_state_0));
    Odrv4 I__699 (
            .O(N__3217),
            .I(my_uart_recv_state_0));
    Odrv4 I__698 (
            .O(N__3214),
            .I(my_uart_recv_state_0));
    LocalMux I__697 (
            .O(N__3209),
            .I(my_uart_recv_state_0));
    InMux I__696 (
            .O(N__3190),
            .I(N__3182));
    InMux I__695 (
            .O(N__3189),
            .I(N__3179));
    InMux I__694 (
            .O(N__3188),
            .I(N__3175));
    InMux I__693 (
            .O(N__3187),
            .I(N__3172));
    InMux I__692 (
            .O(N__3186),
            .I(N__3169));
    InMux I__691 (
            .O(N__3185),
            .I(N__3166));
    LocalMux I__690 (
            .O(N__3182),
            .I(N__3163));
    LocalMux I__689 (
            .O(N__3179),
            .I(N__3160));
    InMux I__688 (
            .O(N__3178),
            .I(N__3157));
    LocalMux I__687 (
            .O(N__3175),
            .I(\my_uart.rx_countdown_3_s1_2 ));
    LocalMux I__686 (
            .O(N__3172),
            .I(\my_uart.rx_countdown_3_s1_2 ));
    LocalMux I__685 (
            .O(N__3169),
            .I(\my_uart.rx_countdown_3_s1_2 ));
    LocalMux I__684 (
            .O(N__3166),
            .I(\my_uart.rx_countdown_3_s1_2 ));
    Odrv12 I__683 (
            .O(N__3163),
            .I(\my_uart.rx_countdown_3_s1_2 ));
    Odrv12 I__682 (
            .O(N__3160),
            .I(\my_uart.rx_countdown_3_s1_2 ));
    LocalMux I__681 (
            .O(N__3157),
            .I(\my_uart.rx_countdown_3_s1_2 ));
    CascadeMux I__680 (
            .O(N__3142),
            .I(N__3139));
    InMux I__679 (
            .O(N__3139),
            .I(N__3136));
    LocalMux I__678 (
            .O(N__3136),
            .I(\my_uart.g0_6_a5_0_4 ));
    InMux I__677 (
            .O(N__3133),
            .I(N__3125));
    InMux I__676 (
            .O(N__3132),
            .I(N__3125));
    InMux I__675 (
            .O(N__3131),
            .I(N__3119));
    InMux I__674 (
            .O(N__3130),
            .I(N__3116));
    LocalMux I__673 (
            .O(N__3125),
            .I(N__3113));
    InMux I__672 (
            .O(N__3124),
            .I(N__3110));
    InMux I__671 (
            .O(N__3123),
            .I(N__3107));
    InMux I__670 (
            .O(N__3122),
            .I(N__3104));
    LocalMux I__669 (
            .O(N__3119),
            .I(\my_uart.rx_countdown_3_s1_4 ));
    LocalMux I__668 (
            .O(N__3116),
            .I(\my_uart.rx_countdown_3_s1_4 ));
    Odrv12 I__667 (
            .O(N__3113),
            .I(\my_uart.rx_countdown_3_s1_4 ));
    LocalMux I__666 (
            .O(N__3110),
            .I(\my_uart.rx_countdown_3_s1_4 ));
    LocalMux I__665 (
            .O(N__3107),
            .I(\my_uart.rx_countdown_3_s1_4 ));
    LocalMux I__664 (
            .O(N__3104),
            .I(\my_uart.rx_countdown_3_s1_4 ));
    InMux I__663 (
            .O(N__3091),
            .I(N__3083));
    InMux I__662 (
            .O(N__3090),
            .I(N__3083));
    InMux I__661 (
            .O(N__3089),
            .I(N__3076));
    InMux I__660 (
            .O(N__3088),
            .I(N__3073));
    LocalMux I__659 (
            .O(N__3083),
            .I(N__3070));
    InMux I__658 (
            .O(N__3082),
            .I(N__3067));
    InMux I__657 (
            .O(N__3081),
            .I(N__3062));
    InMux I__656 (
            .O(N__3080),
            .I(N__3062));
    InMux I__655 (
            .O(N__3079),
            .I(N__3059));
    LocalMux I__654 (
            .O(N__3076),
            .I(\my_uart.rx_countdown_3_s1_5 ));
    LocalMux I__653 (
            .O(N__3073),
            .I(\my_uart.rx_countdown_3_s1_5 ));
    Odrv12 I__652 (
            .O(N__3070),
            .I(\my_uart.rx_countdown_3_s1_5 ));
    LocalMux I__651 (
            .O(N__3067),
            .I(\my_uart.rx_countdown_3_s1_5 ));
    LocalMux I__650 (
            .O(N__3062),
            .I(\my_uart.rx_countdown_3_s1_5 ));
    LocalMux I__649 (
            .O(N__3059),
            .I(\my_uart.rx_countdown_3_s1_5 ));
    InMux I__648 (
            .O(N__3046),
            .I(N__3043));
    LocalMux I__647 (
            .O(N__3043),
            .I(\my_uart.g0_6_a5_0_3 ));
    CascadeMux I__646 (
            .O(N__3040),
            .I(N__3037));
    InMux I__645 (
            .O(N__3037),
            .I(N__3028));
    InMux I__644 (
            .O(N__3036),
            .I(N__3028));
    InMux I__643 (
            .O(N__3035),
            .I(N__3028));
    LocalMux I__642 (
            .O(N__3028),
            .I(\my_uart.rx_bits_remainingZ0Z_1 ));
    InMux I__641 (
            .O(N__3025),
            .I(N__3013));
    InMux I__640 (
            .O(N__3024),
            .I(N__3013));
    InMux I__639 (
            .O(N__3023),
            .I(N__3013));
    InMux I__638 (
            .O(N__3022),
            .I(N__3013));
    LocalMux I__637 (
            .O(N__3013),
            .I(\my_uart.rx_bits_remainingZ0Z_0 ));
    InMux I__636 (
            .O(N__3010),
            .I(N__3007));
    LocalMux I__635 (
            .O(N__3007),
            .I(N__3004));
    Odrv12 I__634 (
            .O(N__3004),
            .I(\my_uart.CO1_i ));
    CascadeMux I__633 (
            .O(N__3001),
            .I(\my_uart.CO1_i_cascade_ ));
    InMux I__632 (
            .O(N__2998),
            .I(N__2995));
    LocalMux I__631 (
            .O(N__2995),
            .I(N__2990));
    InMux I__630 (
            .O(N__2994),
            .I(N__2985));
    InMux I__629 (
            .O(N__2993),
            .I(N__2985));
    Odrv12 I__628 (
            .O(N__2990),
            .I(\my_uart.rx_bits_remainingZ0Z_2 ));
    LocalMux I__627 (
            .O(N__2985),
            .I(\my_uart.rx_bits_remainingZ0Z_2 ));
    CEMux I__626 (
            .O(N__2980),
            .I(N__2977));
    LocalMux I__625 (
            .O(N__2977),
            .I(N__2974));
    Odrv4 I__624 (
            .O(N__2974),
            .I(\my_uart.un1_rx_data_0_sqmuxa_i_i ));
    ClkMux I__623 (
            .O(N__2971),
            .I(N__2932));
    ClkMux I__622 (
            .O(N__2970),
            .I(N__2932));
    ClkMux I__621 (
            .O(N__2969),
            .I(N__2932));
    ClkMux I__620 (
            .O(N__2968),
            .I(N__2932));
    ClkMux I__619 (
            .O(N__2967),
            .I(N__2932));
    ClkMux I__618 (
            .O(N__2966),
            .I(N__2932));
    ClkMux I__617 (
            .O(N__2965),
            .I(N__2932));
    ClkMux I__616 (
            .O(N__2964),
            .I(N__2932));
    ClkMux I__615 (
            .O(N__2963),
            .I(N__2932));
    ClkMux I__614 (
            .O(N__2962),
            .I(N__2932));
    ClkMux I__613 (
            .O(N__2961),
            .I(N__2932));
    ClkMux I__612 (
            .O(N__2960),
            .I(N__2932));
    ClkMux I__611 (
            .O(N__2959),
            .I(N__2932));
    GlobalMux I__610 (
            .O(N__2932),
            .I(N__2929));
    gio2CtrlBuf I__609 (
            .O(N__2929),
            .I(CLK_i_c_g));
    CascadeMux I__608 (
            .O(N__2926),
            .I(\my_uart.m15_e_0_cascade_ ));
    CascadeMux I__607 (
            .O(N__2923),
            .I(\my_uart.m15_e_3_cascade_ ));
    InMux I__606 (
            .O(N__2920),
            .I(N__2917));
    LocalMux I__605 (
            .O(N__2917),
            .I(\my_uart.N_28_mux ));
    InMux I__604 (
            .O(N__2914),
            .I(N__2911));
    LocalMux I__603 (
            .O(N__2911),
            .I(\my_uart.N_19_mux_0 ));
    InMux I__602 (
            .O(N__2908),
            .I(N__2905));
    LocalMux I__601 (
            .O(N__2905),
            .I(\my_uart.m10_e_3 ));
    CascadeMux I__600 (
            .O(N__2902),
            .I(\my_uart.N_19_mux_0_cascade_ ));
    InMux I__599 (
            .O(N__2899),
            .I(N__2892));
    InMux I__598 (
            .O(N__2898),
            .I(N__2882));
    CascadeMux I__597 (
            .O(N__2897),
            .I(N__2878));
    InMux I__596 (
            .O(N__2896),
            .I(N__2872));
    InMux I__595 (
            .O(N__2895),
            .I(N__2872));
    LocalMux I__594 (
            .O(N__2892),
            .I(N__2868));
    InMux I__593 (
            .O(N__2891),
            .I(N__2865));
    CascadeMux I__592 (
            .O(N__2890),
            .I(N__2859));
    InMux I__591 (
            .O(N__2889),
            .I(N__2851));
    InMux I__590 (
            .O(N__2888),
            .I(N__2851));
    InMux I__589 (
            .O(N__2887),
            .I(N__2851));
    InMux I__588 (
            .O(N__2886),
            .I(N__2848));
    InMux I__587 (
            .O(N__2885),
            .I(N__2845));
    LocalMux I__586 (
            .O(N__2882),
            .I(N__2842));
    InMux I__585 (
            .O(N__2881),
            .I(N__2839));
    InMux I__584 (
            .O(N__2878),
            .I(N__2834));
    InMux I__583 (
            .O(N__2877),
            .I(N__2834));
    LocalMux I__582 (
            .O(N__2872),
            .I(N__2831));
    InMux I__581 (
            .O(N__2871),
            .I(N__2828));
    Span4Mux_v I__580 (
            .O(N__2868),
            .I(N__2823));
    LocalMux I__579 (
            .O(N__2865),
            .I(N__2823));
    InMux I__578 (
            .O(N__2864),
            .I(N__2818));
    InMux I__577 (
            .O(N__2863),
            .I(N__2818));
    InMux I__576 (
            .O(N__2862),
            .I(N__2811));
    InMux I__575 (
            .O(N__2859),
            .I(N__2811));
    InMux I__574 (
            .O(N__2858),
            .I(N__2811));
    LocalMux I__573 (
            .O(N__2851),
            .I(\my_uart.un1_rx_clk_divider_a ));
    LocalMux I__572 (
            .O(N__2848),
            .I(\my_uart.un1_rx_clk_divider_a ));
    LocalMux I__571 (
            .O(N__2845),
            .I(\my_uart.un1_rx_clk_divider_a ));
    Odrv4 I__570 (
            .O(N__2842),
            .I(\my_uart.un1_rx_clk_divider_a ));
    LocalMux I__569 (
            .O(N__2839),
            .I(\my_uart.un1_rx_clk_divider_a ));
    LocalMux I__568 (
            .O(N__2834),
            .I(\my_uart.un1_rx_clk_divider_a ));
    Odrv4 I__567 (
            .O(N__2831),
            .I(\my_uart.un1_rx_clk_divider_a ));
    LocalMux I__566 (
            .O(N__2828),
            .I(\my_uart.un1_rx_clk_divider_a ));
    Odrv4 I__565 (
            .O(N__2823),
            .I(\my_uart.un1_rx_clk_divider_a ));
    LocalMux I__564 (
            .O(N__2818),
            .I(\my_uart.un1_rx_clk_divider_a ));
    LocalMux I__563 (
            .O(N__2811),
            .I(\my_uart.un1_rx_clk_divider_a ));
    InMux I__562 (
            .O(N__2788),
            .I(N__2785));
    LocalMux I__561 (
            .O(N__2785),
            .I(\my_uart.N_27_mux ));
    InMux I__560 (
            .O(N__2782),
            .I(N__2773));
    CascadeMux I__559 (
            .O(N__2781),
            .I(N__2769));
    InMux I__558 (
            .O(N__2780),
            .I(N__2763));
    InMux I__557 (
            .O(N__2779),
            .I(N__2763));
    InMux I__556 (
            .O(N__2778),
            .I(N__2760));
    InMux I__555 (
            .O(N__2777),
            .I(N__2757));
    InMux I__554 (
            .O(N__2776),
            .I(N__2754));
    LocalMux I__553 (
            .O(N__2773),
            .I(N__2751));
    InMux I__552 (
            .O(N__2772),
            .I(N__2748));
    InMux I__551 (
            .O(N__2769),
            .I(N__2743));
    InMux I__550 (
            .O(N__2768),
            .I(N__2743));
    LocalMux I__549 (
            .O(N__2763),
            .I(N__2736));
    LocalMux I__548 (
            .O(N__2760),
            .I(N__2736));
    LocalMux I__547 (
            .O(N__2757),
            .I(N__2736));
    LocalMux I__546 (
            .O(N__2754),
            .I(\my_uart.rx_countdownZ0Z_5 ));
    Odrv4 I__545 (
            .O(N__2751),
            .I(\my_uart.rx_countdownZ0Z_5 ));
    LocalMux I__544 (
            .O(N__2748),
            .I(\my_uart.rx_countdownZ0Z_5 ));
    LocalMux I__543 (
            .O(N__2743),
            .I(\my_uart.rx_countdownZ0Z_5 ));
    Odrv4 I__542 (
            .O(N__2736),
            .I(\my_uart.rx_countdownZ0Z_5 ));
    InMux I__541 (
            .O(N__2725),
            .I(N__2722));
    LocalMux I__540 (
            .O(N__2722),
            .I(\my_uart.N_22_mux ));
    CascadeMux I__539 (
            .O(N__2719),
            .I(\my_uart.N_23_mux_cascade_ ));
    InMux I__538 (
            .O(N__2716),
            .I(N__2713));
    LocalMux I__537 (
            .O(N__2713),
            .I(\my_uart.m7_0_0 ));
    InMux I__536 (
            .O(N__2710),
            .I(N__2707));
    LocalMux I__535 (
            .O(N__2707),
            .I(\my_uart.g0_6_0_1 ));
    CascadeMux I__534 (
            .O(N__2704),
            .I(\my_uart.un1_rx_clk_divider28_i_cascade_ ));
    CascadeMux I__533 (
            .O(N__2701),
            .I(N__2693));
    CascadeMux I__532 (
            .O(N__2700),
            .I(N__2690));
    CascadeMux I__531 (
            .O(N__2699),
            .I(N__2682));
    CascadeMux I__530 (
            .O(N__2698),
            .I(N__2678));
    SRMux I__529 (
            .O(N__2697),
            .I(N__2673));
    InMux I__528 (
            .O(N__2696),
            .I(N__2662));
    InMux I__527 (
            .O(N__2693),
            .I(N__2662));
    InMux I__526 (
            .O(N__2690),
            .I(N__2662));
    InMux I__525 (
            .O(N__2689),
            .I(N__2662));
    InMux I__524 (
            .O(N__2688),
            .I(N__2662));
    InMux I__523 (
            .O(N__2687),
            .I(N__2653));
    InMux I__522 (
            .O(N__2686),
            .I(N__2653));
    InMux I__521 (
            .O(N__2685),
            .I(N__2653));
    InMux I__520 (
            .O(N__2682),
            .I(N__2653));
    InMux I__519 (
            .O(N__2681),
            .I(N__2650));
    InMux I__518 (
            .O(N__2678),
            .I(N__2645));
    InMux I__517 (
            .O(N__2677),
            .I(N__2645));
    CascadeMux I__516 (
            .O(N__2676),
            .I(N__2642));
    LocalMux I__515 (
            .O(N__2673),
            .I(N__2637));
    LocalMux I__514 (
            .O(N__2662),
            .I(N__2637));
    LocalMux I__513 (
            .O(N__2653),
            .I(N__2634));
    LocalMux I__512 (
            .O(N__2650),
            .I(N__2627));
    LocalMux I__511 (
            .O(N__2645),
            .I(N__2627));
    InMux I__510 (
            .O(N__2642),
            .I(N__2624));
    Span4Mux_v I__509 (
            .O(N__2637),
            .I(N__2621));
    Span4Mux_h I__508 (
            .O(N__2634),
            .I(N__2618));
    InMux I__507 (
            .O(N__2633),
            .I(N__2613));
    InMux I__506 (
            .O(N__2632),
            .I(N__2613));
    Span4Mux_h I__505 (
            .O(N__2627),
            .I(N__2608));
    LocalMux I__504 (
            .O(N__2624),
            .I(N__2608));
    Odrv4 I__503 (
            .O(N__2621),
            .I(\my_uart.rx_clk_divider_0_sqmuxa ));
    Odrv4 I__502 (
            .O(N__2618),
            .I(\my_uart.rx_clk_divider_0_sqmuxa ));
    LocalMux I__501 (
            .O(N__2613),
            .I(\my_uart.rx_clk_divider_0_sqmuxa ));
    Odrv4 I__500 (
            .O(N__2608),
            .I(\my_uart.rx_clk_divider_0_sqmuxa ));
    InMux I__499 (
            .O(N__2599),
            .I(N__2596));
    LocalMux I__498 (
            .O(N__2596),
            .I(\my_uart.m6_0_18_0 ));
    CascadeMux I__497 (
            .O(N__2593),
            .I(N__2589));
    CascadeMux I__496 (
            .O(N__2592),
            .I(N__2585));
    InMux I__495 (
            .O(N__2589),
            .I(N__2582));
    InMux I__494 (
            .O(N__2588),
            .I(N__2577));
    InMux I__493 (
            .O(N__2585),
            .I(N__2577));
    LocalMux I__492 (
            .O(N__2582),
            .I(N__2574));
    LocalMux I__491 (
            .O(N__2577),
            .I(N__2571));
    Span4Mux_h I__490 (
            .O(N__2574),
            .I(N__2568));
    Odrv4 I__489 (
            .O(N__2571),
            .I(\my_uart.rx_bits_remainingZ0Z_3 ));
    Odrv4 I__488 (
            .O(N__2568),
            .I(\my_uart.rx_bits_remainingZ0Z_3 ));
    InMux I__487 (
            .O(N__2563),
            .I(\my_uart.rx_countdown_3_cry_3_s1 ));
    InMux I__486 (
            .O(N__2560),
            .I(\my_uart.rx_countdown_3_cry_4_s1 ));
    CascadeMux I__485 (
            .O(N__2557),
            .I(N__2554));
    InMux I__484 (
            .O(N__2554),
            .I(N__2547));
    InMux I__483 (
            .O(N__2553),
            .I(N__2547));
    InMux I__482 (
            .O(N__2552),
            .I(N__2544));
    LocalMux I__481 (
            .O(N__2547),
            .I(N__2539));
    LocalMux I__480 (
            .O(N__2544),
            .I(N__2539));
    Span4Mux_v I__479 (
            .O(N__2539),
            .I(N__2534));
    InMux I__478 (
            .O(N__2538),
            .I(N__2531));
    InMux I__477 (
            .O(N__2537),
            .I(N__2528));
    Odrv4 I__476 (
            .O(N__2534),
            .I(\my_uart.un1_recv_state_8 ));
    LocalMux I__475 (
            .O(N__2531),
            .I(\my_uart.un1_recv_state_8 ));
    LocalMux I__474 (
            .O(N__2528),
            .I(\my_uart.un1_recv_state_8 ));
    InMux I__473 (
            .O(N__2521),
            .I(N__2518));
    LocalMux I__472 (
            .O(N__2518),
            .I(N__2515));
    Span4Mux_h I__471 (
            .O(N__2515),
            .I(N__2512));
    Odrv4 I__470 (
            .O(N__2512),
            .I(\my_uart.g0_0_0_a3_3_0 ));
    CascadeMux I__469 (
            .O(N__2509),
            .I(\my_uart.N_8_0_cascade_ ));
    CascadeMux I__468 (
            .O(N__2506),
            .I(N__2503));
    InMux I__467 (
            .O(N__2503),
            .I(N__2500));
    LocalMux I__466 (
            .O(N__2500),
            .I(\my_uart.N_18_mux ));
    CascadeMux I__465 (
            .O(N__2497),
            .I(N__2493));
    CascadeMux I__464 (
            .O(N__2496),
            .I(N__2490));
    InMux I__463 (
            .O(N__2493),
            .I(N__2485));
    InMux I__462 (
            .O(N__2490),
            .I(N__2481));
    CascadeMux I__461 (
            .O(N__2489),
            .I(N__2477));
    CascadeMux I__460 (
            .O(N__2488),
            .I(N__2474));
    LocalMux I__459 (
            .O(N__2485),
            .I(N__2471));
    CascadeMux I__458 (
            .O(N__2484),
            .I(N__2466));
    LocalMux I__457 (
            .O(N__2481),
            .I(N__2463));
    InMux I__456 (
            .O(N__2480),
            .I(N__2458));
    InMux I__455 (
            .O(N__2477),
            .I(N__2458));
    InMux I__454 (
            .O(N__2474),
            .I(N__2455));
    Span4Mux_v I__453 (
            .O(N__2471),
            .I(N__2452));
    InMux I__452 (
            .O(N__2470),
            .I(N__2447));
    InMux I__451 (
            .O(N__2469),
            .I(N__2447));
    InMux I__450 (
            .O(N__2466),
            .I(N__2444));
    Odrv4 I__449 (
            .O(N__2463),
            .I(\my_uart.rx_countdownZ0Z_4 ));
    LocalMux I__448 (
            .O(N__2458),
            .I(\my_uart.rx_countdownZ0Z_4 ));
    LocalMux I__447 (
            .O(N__2455),
            .I(\my_uart.rx_countdownZ0Z_4 ));
    Odrv4 I__446 (
            .O(N__2452),
            .I(\my_uart.rx_countdownZ0Z_4 ));
    LocalMux I__445 (
            .O(N__2447),
            .I(\my_uart.rx_countdownZ0Z_4 ));
    LocalMux I__444 (
            .O(N__2444),
            .I(\my_uart.rx_countdownZ0Z_4 ));
    InMux I__443 (
            .O(N__2431),
            .I(N__2428));
    LocalMux I__442 (
            .O(N__2428),
            .I(N__2422));
    CascadeMux I__441 (
            .O(N__2427),
            .I(N__2414));
    InMux I__440 (
            .O(N__2426),
            .I(N__2409));
    InMux I__439 (
            .O(N__2425),
            .I(N__2409));
    Span4Mux_v I__438 (
            .O(N__2422),
            .I(N__2406));
    InMux I__437 (
            .O(N__2421),
            .I(N__2403));
    InMux I__436 (
            .O(N__2420),
            .I(N__2400));
    InMux I__435 (
            .O(N__2419),
            .I(N__2397));
    InMux I__434 (
            .O(N__2418),
            .I(N__2392));
    InMux I__433 (
            .O(N__2417),
            .I(N__2392));
    InMux I__432 (
            .O(N__2414),
            .I(N__2389));
    LocalMux I__431 (
            .O(N__2409),
            .I(\my_uart.rx_countdownZ1Z_1 ));
    Odrv4 I__430 (
            .O(N__2406),
            .I(\my_uart.rx_countdownZ1Z_1 ));
    LocalMux I__429 (
            .O(N__2403),
            .I(\my_uart.rx_countdownZ1Z_1 ));
    LocalMux I__428 (
            .O(N__2400),
            .I(\my_uart.rx_countdownZ1Z_1 ));
    LocalMux I__427 (
            .O(N__2397),
            .I(\my_uart.rx_countdownZ1Z_1 ));
    LocalMux I__426 (
            .O(N__2392),
            .I(\my_uart.rx_countdownZ1Z_1 ));
    LocalMux I__425 (
            .O(N__2389),
            .I(\my_uart.rx_countdownZ1Z_1 ));
    InMux I__424 (
            .O(N__2374),
            .I(N__2371));
    LocalMux I__423 (
            .O(N__2371),
            .I(N__2363));
    CascadeMux I__422 (
            .O(N__2370),
            .I(N__2358));
    InMux I__421 (
            .O(N__2369),
            .I(N__2355));
    InMux I__420 (
            .O(N__2368),
            .I(N__2352));
    InMux I__419 (
            .O(N__2367),
            .I(N__2347));
    InMux I__418 (
            .O(N__2366),
            .I(N__2347));
    Span4Mux_h I__417 (
            .O(N__2363),
            .I(N__2344));
    InMux I__416 (
            .O(N__2362),
            .I(N__2339));
    InMux I__415 (
            .O(N__2361),
            .I(N__2339));
    InMux I__414 (
            .O(N__2358),
            .I(N__2336));
    LocalMux I__413 (
            .O(N__2355),
            .I(\my_uart.rx_countdownZ1Z_2 ));
    LocalMux I__412 (
            .O(N__2352),
            .I(\my_uart.rx_countdownZ1Z_2 ));
    LocalMux I__411 (
            .O(N__2347),
            .I(\my_uart.rx_countdownZ1Z_2 ));
    Odrv4 I__410 (
            .O(N__2344),
            .I(\my_uart.rx_countdownZ1Z_2 ));
    LocalMux I__409 (
            .O(N__2339),
            .I(\my_uart.rx_countdownZ1Z_2 ));
    LocalMux I__408 (
            .O(N__2336),
            .I(\my_uart.rx_countdownZ1Z_2 ));
    InMux I__407 (
            .O(N__2323),
            .I(N__2319));
    InMux I__406 (
            .O(N__2322),
            .I(N__2315));
    LocalMux I__405 (
            .O(N__2319),
            .I(N__2309));
    InMux I__404 (
            .O(N__2318),
            .I(N__2306));
    LocalMux I__403 (
            .O(N__2315),
            .I(N__2301));
    InMux I__402 (
            .O(N__2314),
            .I(N__2298));
    InMux I__401 (
            .O(N__2313),
            .I(N__2293));
    InMux I__400 (
            .O(N__2312),
            .I(N__2293));
    Span4Mux_h I__399 (
            .O(N__2309),
            .I(N__2290));
    LocalMux I__398 (
            .O(N__2306),
            .I(N__2287));
    InMux I__397 (
            .O(N__2305),
            .I(N__2284));
    InMux I__396 (
            .O(N__2304),
            .I(N__2281));
    Odrv4 I__395 (
            .O(N__2301),
            .I(\my_uart.rx_countdownZ1Z_3 ));
    LocalMux I__394 (
            .O(N__2298),
            .I(\my_uart.rx_countdownZ1Z_3 ));
    LocalMux I__393 (
            .O(N__2293),
            .I(\my_uart.rx_countdownZ1Z_3 ));
    Odrv4 I__392 (
            .O(N__2290),
            .I(\my_uart.rx_countdownZ1Z_3 ));
    Odrv4 I__391 (
            .O(N__2287),
            .I(\my_uart.rx_countdownZ1Z_3 ));
    LocalMux I__390 (
            .O(N__2284),
            .I(\my_uart.rx_countdownZ1Z_3 ));
    LocalMux I__389 (
            .O(N__2281),
            .I(\my_uart.rx_countdownZ1Z_3 ));
    CascadeMux I__388 (
            .O(N__2266),
            .I(\my_uart.m10_e_1_cascade_ ));
    CascadeMux I__387 (
            .O(N__2263),
            .I(\my_uart.g0_4_a3_3_cascade_ ));
    InMux I__386 (
            .O(N__2260),
            .I(N__2257));
    LocalMux I__385 (
            .O(N__2257),
            .I(\my_uart.g0_4_a3_4 ));
    InMux I__384 (
            .O(N__2254),
            .I(N__2251));
    LocalMux I__383 (
            .O(N__2251),
            .I(\my_uart.recv_state_0_sqmuxa_1_0 ));
    InMux I__382 (
            .O(N__2248),
            .I(N__2245));
    LocalMux I__381 (
            .O(N__2245),
            .I(\my_uart.g0_4_a3_0_2 ));
    InMux I__380 (
            .O(N__2242),
            .I(N__2239));
    LocalMux I__379 (
            .O(N__2239),
            .I(\my_uart.g0_6_a5_1_0 ));
    InMux I__378 (
            .O(N__2236),
            .I(\my_uart.rx_countdown_3_cry_0_s1 ));
    InMux I__377 (
            .O(N__2233),
            .I(\my_uart.rx_countdown_3_cry_1_s1 ));
    InMux I__376 (
            .O(N__2230),
            .I(\my_uart.rx_countdown_3_cry_2_s1 ));
    CascadeMux I__375 (
            .O(N__2227),
            .I(N__2222));
    CascadeMux I__374 (
            .O(N__2226),
            .I(N__2217));
    InMux I__373 (
            .O(N__2225),
            .I(N__2210));
    InMux I__372 (
            .O(N__2222),
            .I(N__2210));
    InMux I__371 (
            .O(N__2221),
            .I(N__2210));
    InMux I__370 (
            .O(N__2220),
            .I(N__2204));
    InMux I__369 (
            .O(N__2217),
            .I(N__2204));
    LocalMux I__368 (
            .O(N__2210),
            .I(N__2194));
    InMux I__367 (
            .O(N__2209),
            .I(N__2191));
    LocalMux I__366 (
            .O(N__2204),
            .I(N__2188));
    CascadeMux I__365 (
            .O(N__2203),
            .I(N__2185));
    CascadeMux I__364 (
            .O(N__2202),
            .I(N__2182));
    CascadeMux I__363 (
            .O(N__2201),
            .I(N__2179));
    CascadeMux I__362 (
            .O(N__2200),
            .I(N__2176));
    CascadeMux I__361 (
            .O(N__2199),
            .I(N__2173));
    CascadeMux I__360 (
            .O(N__2198),
            .I(N__2170));
    CascadeMux I__359 (
            .O(N__2197),
            .I(N__2167));
    Span4Mux_v I__358 (
            .O(N__2194),
            .I(N__2164));
    LocalMux I__357 (
            .O(N__2191),
            .I(N__2161));
    Span4Mux_v I__356 (
            .O(N__2188),
            .I(N__2158));
    InMux I__355 (
            .O(N__2185),
            .I(N__2151));
    InMux I__354 (
            .O(N__2182),
            .I(N__2151));
    InMux I__353 (
            .O(N__2179),
            .I(N__2151));
    InMux I__352 (
            .O(N__2176),
            .I(N__2142));
    InMux I__351 (
            .O(N__2173),
            .I(N__2142));
    InMux I__350 (
            .O(N__2170),
            .I(N__2142));
    InMux I__349 (
            .O(N__2167),
            .I(N__2142));
    Odrv4 I__348 (
            .O(N__2164),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__347 (
            .O(N__2161),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__346 (
            .O(N__2158),
            .I(CONSTANT_ONE_NET));
    LocalMux I__345 (
            .O(N__2151),
            .I(CONSTANT_ONE_NET));
    LocalMux I__344 (
            .O(N__2142),
            .I(CONSTANT_ONE_NET));
    InMux I__343 (
            .O(N__2131),
            .I(N__2128));
    LocalMux I__342 (
            .O(N__2128),
            .I(\my_uart.rx_countdown_3_4 ));
    CascadeMux I__341 (
            .O(N__2125),
            .I(\my_uart.rx_countdown_3_4_cascade_ ));
    InMux I__340 (
            .O(N__2122),
            .I(N__2119));
    LocalMux I__339 (
            .O(N__2119),
            .I(N__2116));
    Odrv4 I__338 (
            .O(N__2116),
            .I(\my_uart.rx_countdown_RNO_4Z0Z_2 ));
    InMux I__337 (
            .O(N__2113),
            .I(N__2110));
    LocalMux I__336 (
            .O(N__2110),
            .I(\my_uart.N_13 ));
    InMux I__335 (
            .O(N__2107),
            .I(N__2101));
    InMux I__334 (
            .O(N__2106),
            .I(N__2101));
    LocalMux I__333 (
            .O(N__2101),
            .I(\my_uart.rx_countdown_3_3 ));
    InMux I__332 (
            .O(N__2098),
            .I(N__2095));
    LocalMux I__331 (
            .O(N__2095),
            .I(\my_uart.G_14_0_a3_0_1 ));
    InMux I__330 (
            .O(N__2092),
            .I(N__2089));
    LocalMux I__329 (
            .O(N__2089),
            .I(\my_uart.g0_6_0_0 ));
    CascadeMux I__328 (
            .O(N__2086),
            .I(N__2083));
    InMux I__327 (
            .O(N__2083),
            .I(N__2080));
    LocalMux I__326 (
            .O(N__2080),
            .I(\my_uart.g0_4_a3_0_3 ));
    CascadeMux I__325 (
            .O(N__2077),
            .I(\my_uart.rx_countdown20_cascade_ ));
    InMux I__324 (
            .O(N__2074),
            .I(N__2071));
    LocalMux I__323 (
            .O(N__2071),
            .I(\my_uart.un1_recv_state_6 ));
    InMux I__322 (
            .O(N__2068),
            .I(N__2065));
    LocalMux I__321 (
            .O(N__2065),
            .I(N__2060));
    InMux I__320 (
            .O(N__2064),
            .I(N__2057));
    CEMux I__319 (
            .O(N__2063),
            .I(N__2054));
    Span4Mux_h I__318 (
            .O(N__2060),
            .I(N__2051));
    LocalMux I__317 (
            .O(N__2057),
            .I(\my_uart.rx_data_0_sqmuxa ));
    LocalMux I__316 (
            .O(N__2054),
            .I(\my_uart.rx_data_0_sqmuxa ));
    Odrv4 I__315 (
            .O(N__2051),
            .I(\my_uart.rx_data_0_sqmuxa ));
    CascadeMux I__314 (
            .O(N__2044),
            .I(\my_uart.N_6_cascade_ ));
    InMux I__313 (
            .O(N__2041),
            .I(N__2038));
    LocalMux I__312 (
            .O(N__2038),
            .I(\my_uart.un1_rx_clk_divider_a_0 ));
    CascadeMux I__311 (
            .O(N__2035),
            .I(N__2030));
    InMux I__310 (
            .O(N__2034),
            .I(N__2027));
    InMux I__309 (
            .O(N__2033),
            .I(N__2024));
    InMux I__308 (
            .O(N__2030),
            .I(N__2021));
    LocalMux I__307 (
            .O(N__2027),
            .I(N__2018));
    LocalMux I__306 (
            .O(N__2024),
            .I(\my_uart.rx_clk_dividerZ0Z_9 ));
    LocalMux I__305 (
            .O(N__2021),
            .I(\my_uart.rx_clk_dividerZ0Z_9 ));
    Odrv4 I__304 (
            .O(N__2018),
            .I(\my_uart.rx_clk_dividerZ0Z_9 ));
    CascadeMux I__303 (
            .O(N__2011),
            .I(N__2008));
    InMux I__302 (
            .O(N__2008),
            .I(N__2005));
    LocalMux I__301 (
            .O(N__2005),
            .I(\my_uart.un1_rx_clk_divider_a_6 ));
    InMux I__300 (
            .O(N__2002),
            .I(N__1999));
    LocalMux I__299 (
            .O(N__1999),
            .I(N__1996));
    Odrv4 I__298 (
            .O(N__1996),
            .I(\my_uart.un1_rx_clk_divider_a_7 ));
    CascadeMux I__297 (
            .O(N__1993),
            .I(\my_uart.un1_rx_clk_divider_a_cascade_ ));
    InMux I__296 (
            .O(N__1990),
            .I(N__1987));
    LocalMux I__295 (
            .O(N__1987),
            .I(N__1984));
    Odrv4 I__294 (
            .O(N__1984),
            .I(\my_uart.N_5 ));
    InMux I__293 (
            .O(N__1981),
            .I(N__1978));
    LocalMux I__292 (
            .O(N__1978),
            .I(\my_uart.g0_0_0_a3_0_3 ));
    CascadeMux I__291 (
            .O(N__1975),
            .I(\my_uart.g0_6_a5_1_5_cascade_ ));
    InMux I__290 (
            .O(N__1972),
            .I(N__1969));
    LocalMux I__289 (
            .O(N__1969),
            .I(\my_uart.g0_6_a5_1_4 ));
    CascadeMux I__288 (
            .O(N__1966),
            .I(\my_uart.rx_countdown_8_5_cascade_ ));
    InMux I__287 (
            .O(N__1963),
            .I(N__1956));
    InMux I__286 (
            .O(N__1962),
            .I(N__1956));
    InMux I__285 (
            .O(N__1961),
            .I(N__1953));
    LocalMux I__284 (
            .O(N__1956),
            .I(\my_uart.rx_clk_dividerZ0Z_8 ));
    LocalMux I__283 (
            .O(N__1953),
            .I(\my_uart.rx_clk_dividerZ0Z_8 ));
    InMux I__282 (
            .O(N__1948),
            .I(N__1945));
    LocalMux I__281 (
            .O(N__1945),
            .I(\my_uart.rx_countdown_RNO_5Z0Z_2 ));
    CascadeMux I__280 (
            .O(N__1942),
            .I(\my_uart.rx_countdown_RNO_6Z0Z_2_cascade_ ));
    InMux I__279 (
            .O(N__1939),
            .I(N__1936));
    LocalMux I__278 (
            .O(N__1936),
            .I(\my_uart.rx_clk_divider_1_cry_6_THRU_CO ));
    InMux I__277 (
            .O(N__1933),
            .I(N__1928));
    InMux I__276 (
            .O(N__1932),
            .I(N__1923));
    InMux I__275 (
            .O(N__1931),
            .I(N__1923));
    LocalMux I__274 (
            .O(N__1928),
            .I(\my_uart.rx_clk_dividerZ0Z_7 ));
    LocalMux I__273 (
            .O(N__1923),
            .I(\my_uart.rx_clk_dividerZ0Z_7 ));
    InMux I__272 (
            .O(N__1918),
            .I(N__1915));
    LocalMux I__271 (
            .O(N__1915),
            .I(\my_uart.rx_clk_divider_1_cry_7_THRU_CO ));
    InMux I__270 (
            .O(N__1912),
            .I(N__1909));
    LocalMux I__269 (
            .O(N__1909),
            .I(\my_uart.rx_clk_divider_1_cry_8_THRU_CO ));
    InMux I__268 (
            .O(N__1906),
            .I(N__1903));
    LocalMux I__267 (
            .O(N__1903),
            .I(\my_uart.rx_clk_divider_1_cry_1_THRU_CO ));
    InMux I__266 (
            .O(N__1900),
            .I(N__1895));
    InMux I__265 (
            .O(N__1899),
            .I(N__1890));
    InMux I__264 (
            .O(N__1898),
            .I(N__1890));
    LocalMux I__263 (
            .O(N__1895),
            .I(\my_uart.rx_clk_dividerZ0Z_2 ));
    LocalMux I__262 (
            .O(N__1890),
            .I(\my_uart.rx_clk_dividerZ0Z_2 ));
    InMux I__261 (
            .O(N__1885),
            .I(N__1882));
    LocalMux I__260 (
            .O(N__1882),
            .I(N__1879));
    Odrv4 I__259 (
            .O(N__1879),
            .I(\my_uart.rx_clk_divider_1_cry_2_THRU_CO ));
    InMux I__258 (
            .O(N__1876),
            .I(N__1873));
    LocalMux I__257 (
            .O(N__1873),
            .I(N__1870));
    Odrv4 I__256 (
            .O(N__1870),
            .I(\my_uart.rx_clk_divider_1_cry_3_THRU_CO ));
    InMux I__255 (
            .O(N__1867),
            .I(N__1864));
    LocalMux I__254 (
            .O(N__1864),
            .I(N__1861));
    Odrv4 I__253 (
            .O(N__1861),
            .I(\my_uart.rx_clk_divider_1_cry_5_THRU_CO ));
    InMux I__252 (
            .O(N__1858),
            .I(N__1855));
    LocalMux I__251 (
            .O(N__1855),
            .I(N__1852));
    Odrv4 I__250 (
            .O(N__1852),
            .I(\my_uart.rx_clk_divider_1_cry_4_THRU_CO ));
    InMux I__249 (
            .O(N__1849),
            .I(N__1845));
    CascadeMux I__248 (
            .O(N__1848),
            .I(N__1842));
    LocalMux I__247 (
            .O(N__1845),
            .I(N__1838));
    InMux I__246 (
            .O(N__1842),
            .I(N__1833));
    InMux I__245 (
            .O(N__1841),
            .I(N__1833));
    Odrv4 I__244 (
            .O(N__1838),
            .I(\my_uart.rx_clk_dividerZ0Z_5 ));
    LocalMux I__243 (
            .O(N__1833),
            .I(\my_uart.rx_clk_dividerZ0Z_5 ));
    CascadeMux I__242 (
            .O(N__1828),
            .I(N__1824));
    InMux I__241 (
            .O(N__1827),
            .I(N__1821));
    InMux I__240 (
            .O(N__1824),
            .I(N__1817));
    LocalMux I__239 (
            .O(N__1821),
            .I(N__1814));
    InMux I__238 (
            .O(N__1820),
            .I(N__1811));
    LocalMux I__237 (
            .O(N__1817),
            .I(\my_uart.rx_clk_dividerZ0Z_4 ));
    Odrv4 I__236 (
            .O(N__1814),
            .I(\my_uart.rx_clk_dividerZ0Z_4 ));
    LocalMux I__235 (
            .O(N__1811),
            .I(\my_uart.rx_clk_dividerZ0Z_4 ));
    InMux I__234 (
            .O(N__1804),
            .I(N__1800));
    CascadeMux I__233 (
            .O(N__1803),
            .I(N__1796));
    LocalMux I__232 (
            .O(N__1800),
            .I(N__1793));
    InMux I__231 (
            .O(N__1799),
            .I(N__1788));
    InMux I__230 (
            .O(N__1796),
            .I(N__1788));
    Odrv4 I__229 (
            .O(N__1793),
            .I(\my_uart.rx_clk_dividerZ0Z_6 ));
    LocalMux I__228 (
            .O(N__1788),
            .I(\my_uart.rx_clk_dividerZ0Z_6 ));
    InMux I__227 (
            .O(N__1783),
            .I(N__1780));
    LocalMux I__226 (
            .O(N__1780),
            .I(N__1775));
    InMux I__225 (
            .O(N__1779),
            .I(N__1770));
    InMux I__224 (
            .O(N__1778),
            .I(N__1770));
    Odrv4 I__223 (
            .O(N__1775),
            .I(\my_uart.rx_clk_dividerZ0Z_3 ));
    LocalMux I__222 (
            .O(N__1770),
            .I(\my_uart.rx_clk_dividerZ0Z_3 ));
    InMux I__221 (
            .O(N__1765),
            .I(\my_uart.rx_clk_divider_1_cry_3 ));
    InMux I__220 (
            .O(N__1762),
            .I(\my_uart.rx_clk_divider_1_cry_4 ));
    InMux I__219 (
            .O(N__1759),
            .I(\my_uart.rx_clk_divider_1_cry_5 ));
    InMux I__218 (
            .O(N__1756),
            .I(\my_uart.rx_clk_divider_1_cry_6 ));
    InMux I__217 (
            .O(N__1753),
            .I(bfn_9_26_0_));
    InMux I__216 (
            .O(N__1750),
            .I(\my_uart.rx_clk_divider_1_cry_8 ));
    InMux I__215 (
            .O(N__1747),
            .I(\my_uart.rx_clk_divider_1_cry_9 ));
    InMux I__214 (
            .O(N__1744),
            .I(N__1740));
    InMux I__213 (
            .O(N__1743),
            .I(N__1737));
    LocalMux I__212 (
            .O(N__1740),
            .I(\my_uart.rx_clk_dividerZ0Z_1 ));
    LocalMux I__211 (
            .O(N__1737),
            .I(\my_uart.rx_clk_dividerZ0Z_1 ));
    CascadeMux I__210 (
            .O(N__1732),
            .I(N__1728));
    InMux I__209 (
            .O(N__1731),
            .I(N__1725));
    InMux I__208 (
            .O(N__1728),
            .I(N__1722));
    LocalMux I__207 (
            .O(N__1725),
            .I(\my_uart.rx_clk_dividerZ0Z_10 ));
    LocalMux I__206 (
            .O(N__1722),
            .I(\my_uart.rx_clk_dividerZ0Z_10 ));
    InMux I__205 (
            .O(N__1717),
            .I(N__1714));
    LocalMux I__204 (
            .O(N__1714),
            .I(\my_uart.rx_clk_divider_1_cry_0_THRU_CO ));
    InMux I__203 (
            .O(N__1711),
            .I(N__1706));
    InMux I__202 (
            .O(N__1710),
            .I(N__1701));
    InMux I__201 (
            .O(N__1709),
            .I(N__1701));
    LocalMux I__200 (
            .O(N__1706),
            .I(\my_uart.rx_clk_dividerZ1Z_1 ));
    LocalMux I__199 (
            .O(N__1701),
            .I(\my_uart.rx_clk_dividerZ1Z_1 ));
    IoInMux I__198 (
            .O(N__1696),
            .I(N__1693));
    LocalMux I__197 (
            .O(N__1693),
            .I(N__1690));
    IoSpan4Mux I__196 (
            .O(N__1690),
            .I(N__1687));
    Span4Mux_s1_v I__195 (
            .O(N__1687),
            .I(N__1684));
    Span4Mux_v I__194 (
            .O(N__1684),
            .I(N__1680));
    InMux I__193 (
            .O(N__1683),
            .I(N__1677));
    Odrv4 I__192 (
            .O(N__1680),
            .I(LED_o_c_7));
    LocalMux I__191 (
            .O(N__1677),
            .I(LED_o_c_7));
    IoInMux I__190 (
            .O(N__1672),
            .I(N__1669));
    LocalMux I__189 (
            .O(N__1669),
            .I(N__1666));
    Span4Mux_s2_v I__188 (
            .O(N__1666),
            .I(N__1663));
    Span4Mux_h I__187 (
            .O(N__1663),
            .I(N__1659));
    InMux I__186 (
            .O(N__1662),
            .I(N__1656));
    Odrv4 I__185 (
            .O(N__1659),
            .I(LED_o_c_6));
    LocalMux I__184 (
            .O(N__1656),
            .I(LED_o_c_6));
    IoInMux I__183 (
            .O(N__1651),
            .I(N__1648));
    LocalMux I__182 (
            .O(N__1648),
            .I(N__1645));
    IoSpan4Mux I__181 (
            .O(N__1645),
            .I(N__1642));
    Span4Mux_s2_v I__180 (
            .O(N__1642),
            .I(N__1638));
    InMux I__179 (
            .O(N__1641),
            .I(N__1635));
    Odrv4 I__178 (
            .O(N__1638),
            .I(LED_o_c_3));
    LocalMux I__177 (
            .O(N__1635),
            .I(LED_o_c_3));
    IoInMux I__176 (
            .O(N__1630),
            .I(N__1627));
    LocalMux I__175 (
            .O(N__1627),
            .I(N__1624));
    IoSpan4Mux I__174 (
            .O(N__1624),
            .I(N__1621));
    Span4Mux_s2_v I__173 (
            .O(N__1621),
            .I(N__1617));
    InMux I__172 (
            .O(N__1620),
            .I(N__1614));
    Odrv4 I__171 (
            .O(N__1617),
            .I(LED_o_c_2));
    LocalMux I__170 (
            .O(N__1614),
            .I(LED_o_c_2));
    IoInMux I__169 (
            .O(N__1609),
            .I(N__1606));
    LocalMux I__168 (
            .O(N__1606),
            .I(N__1603));
    Span4Mux_s1_v I__167 (
            .O(N__1603),
            .I(N__1600));
    Span4Mux_v I__166 (
            .O(N__1600),
            .I(N__1596));
    InMux I__165 (
            .O(N__1599),
            .I(N__1593));
    Odrv4 I__164 (
            .O(N__1596),
            .I(LED_o_c_1));
    LocalMux I__163 (
            .O(N__1593),
            .I(LED_o_c_1));
    IoInMux I__162 (
            .O(N__1588),
            .I(N__1585));
    LocalMux I__161 (
            .O(N__1585),
            .I(N__1582));
    Span4Mux_s2_v I__160 (
            .O(N__1582),
            .I(N__1579));
    Span4Mux_h I__159 (
            .O(N__1579),
            .I(N__1575));
    InMux I__158 (
            .O(N__1578),
            .I(N__1572));
    Odrv4 I__157 (
            .O(N__1575),
            .I(LED_o_c_5));
    LocalMux I__156 (
            .O(N__1572),
            .I(LED_o_c_5));
    IoInMux I__155 (
            .O(N__1567),
            .I(N__1564));
    LocalMux I__154 (
            .O(N__1564),
            .I(N__1561));
    Span12Mux_s5_v I__153 (
            .O(N__1561),
            .I(N__1557));
    InMux I__152 (
            .O(N__1560),
            .I(N__1554));
    Odrv12 I__151 (
            .O(N__1557),
            .I(LED_o_c_4));
    LocalMux I__150 (
            .O(N__1554),
            .I(LED_o_c_4));
    InMux I__149 (
            .O(N__1549),
            .I(\my_uart.rx_clk_divider_1_cry_0 ));
    InMux I__148 (
            .O(N__1546),
            .I(\my_uart.rx_clk_divider_1_cry_1 ));
    InMux I__147 (
            .O(N__1543),
            .I(\my_uart.rx_clk_divider_1_cry_2 ));
    InMux I__146 (
            .O(N__1540),
            .I(N__1537));
    LocalMux I__145 (
            .O(N__1537),
            .I(\my_uart.rx_bits_remaining_6_0_3 ));
    CascadeMux I__144 (
            .O(N__1534),
            .I(\my_uart.g0_0_0_a3_3_cascade_ ));
    CascadeMux I__143 (
            .O(N__1531),
            .I(\my_uart.N_4_cascade_ ));
    InMux I__142 (
            .O(N__1528),
            .I(N__1525));
    LocalMux I__141 (
            .O(N__1525),
            .I(N__1522));
    Odrv4 I__140 (
            .O(N__1522),
            .I(\my_uart.g0_0 ));
    InMux I__139 (
            .O(N__1519),
            .I(N__1516));
    LocalMux I__138 (
            .O(N__1516),
            .I(\my_uart.g0_0_0_a3_4 ));
    IoInMux I__137 (
            .O(N__1513),
            .I(N__1510));
    LocalMux I__136 (
            .O(N__1510),
            .I(N__1507));
    Odrv12 I__135 (
            .O(N__1507),
            .I(LED_o_c_0));
    CascadeMux I__134 (
            .O(N__1504),
            .I(\my_uart.recv_state_0_sqmuxa_1_cascade_ ));
    CascadeMux I__133 (
            .O(N__1501),
            .I(N__1498));
    InMux I__132 (
            .O(N__1498),
            .I(N__1495));
    LocalMux I__131 (
            .O(N__1495),
            .I(N__1492));
    Odrv4 I__130 (
            .O(N__1492),
            .I(\my_uart.g0_2 ));
    CascadeMux I__129 (
            .O(N__1489),
            .I(\my_uart.g0_0_0_a3_0_0_cascade_ ));
    InMux I__128 (
            .O(N__1486),
            .I(N__1483));
    LocalMux I__127 (
            .O(N__1483),
            .I(\my_uart.g0_0_0_a3_0_4 ));
    defparam IN_MUX_bfv_9_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_25_0_));
    defparam IN_MUX_bfv_9_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_26_0_ (
            .carryinitin(\my_uart.rx_clk_divider_1_cry_7 ),
            .carryinitout(bfn_9_26_0_));
    defparam IN_MUX_bfv_11_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_26_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \my_uart.rx_bits_remaining_RNO_0_3_LC_7_25_0 .C_ON=1'b0;
    defparam \my_uart.rx_bits_remaining_RNO_0_3_LC_7_25_0 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_bits_remaining_RNO_0_3_LC_7_25_0 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \my_uart.rx_bits_remaining_RNO_0_3_LC_7_25_0  (
            .in0(N__1486),
            .in1(N__2899),
            .in2(N__1501),
            .in3(N__1519),
            .lcout(),
            .ltout(\my_uart.recv_state_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_bits_remaining_3_LC_7_25_1 .C_ON=1'b0;
    defparam \my_uart.rx_bits_remaining_3_LC_7_25_1 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_bits_remaining_3_LC_7_25_1 .LUT_INIT=16'b0011001100111010;
    LogicCell40 \my_uart.rx_bits_remaining_3_LC_7_25_1  (
            .in0(N__2588),
            .in1(N__1540),
            .in2(N__1504),
            .in3(N__2064),
            .lcout(\my_uart.rx_bits_remainingZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2959),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_bits_remaining_RNO_4_3_LC_7_25_4 .C_ON=1'b0;
    defparam \my_uart.rx_bits_remaining_RNO_4_3_LC_7_25_4 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_bits_remaining_RNO_4_3_LC_7_25_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \my_uart.rx_bits_remaining_RNO_4_3_LC_7_25_4  (
            .in0(N__3567),
            .in1(N__3305),
            .in2(N__3841),
            .in3(N__3454),
            .lcout(\my_uart.g0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_bits_remaining_RNO_5_3_LC_7_25_5 .C_ON=1'b0;
    defparam \my_uart.rx_bits_remaining_RNO_5_3_LC_7_25_5 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_bits_remaining_RNO_5_3_LC_7_25_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \my_uart.rx_bits_remaining_RNO_5_3_LC_7_25_5  (
            .in0(N__2323),
            .in1(N__2374),
            .in2(N__2497),
            .in3(N__3667),
            .lcout(),
            .ltout(\my_uart.g0_0_0_a3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_bits_remaining_RNO_2_3_LC_7_25_6 .C_ON=1'b0;
    defparam \my_uart.rx_bits_remaining_RNO_2_3_LC_7_25_6 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_bits_remaining_RNO_2_3_LC_7_25_6 .LUT_INIT=16'b0001000000010000;
    LogicCell40 \my_uart.rx_bits_remaining_RNO_2_3_LC_7_25_6  (
            .in0(N__2431),
            .in1(N__2782),
            .in2(N__1489),
            .in3(_gnd_net_),
            .lcout(\my_uart.g0_0_0_a3_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_bits_remaining_RNO_1_3_LC_7_25_7 .C_ON=1'b0;
    defparam \my_uart.rx_bits_remaining_RNO_1_3_LC_7_25_7 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_bits_remaining_RNO_1_3_LC_7_25_7 .LUT_INIT=16'b0001010000000101;
    LogicCell40 \my_uart.rx_bits_remaining_RNO_1_3_LC_7_25_7  (
            .in0(N__3306),
            .in1(N__2998),
            .in2(N__2592),
            .in3(N__3010),
            .lcout(\my_uart.rx_bits_remaining_6_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_RNIH36N1_0_LC_7_26_0 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_RNIH36N1_0_LC_7_26_0 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_RNIH36N1_0_LC_7_26_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \my_uart.rx_countdown_RNIH36N1_0_LC_7_26_0  (
            .in0(N__3190),
            .in1(N__3666),
            .in2(N__3367),
            .in3(N__3718),
            .lcout(),
            .ltout(\my_uart.g0_0_0_a3_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_RNIPOKB5_0_LC_7_26_1 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_RNIPOKB5_0_LC_7_26_1 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_RNIPOKB5_0_LC_7_26_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \my_uart.rx_countdown_RNIPOKB5_0_LC_7_26_1  (
            .in0(N__3091),
            .in1(N__3133),
            .in2(N__1534),
            .in3(N__2891),
            .lcout(),
            .ltout(\my_uart.N_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNI4O0M9_2_LC_7_26_2 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNI4O0M9_2_LC_7_26_2 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNI4O0M9_2_LC_7_26_2 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \my_uart.recv_state_RNI4O0M9_2_LC_7_26_2  (
            .in0(N__1990),
            .in1(N__3568),
            .in2(N__1531),
            .in3(N__1528),
            .lcout(\my_uart.rx_data_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNIF559_1_LC_7_26_4 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNIF559_1_LC_7_26_4 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNIF559_1_LC_7_26_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \my_uart.recv_state_RNIF559_1_LC_7_26_4  (
            .in0(_gnd_net_),
            .in1(N__3310),
            .in2(_gnd_net_),
            .in3(N__3460),
            .lcout(\my_uart.g0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_bits_remaining_RNO_3_3_LC_7_26_5 .C_ON=1'b0;
    defparam \my_uart.rx_bits_remaining_RNO_3_3_LC_7_26_5 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_bits_remaining_RNO_3_3_LC_7_26_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \my_uart.rx_bits_remaining_RNO_3_3_LC_7_26_5  (
            .in0(N__3090),
            .in1(N__3132),
            .in2(_gnd_net_),
            .in3(N__2521),
            .lcout(\my_uart.g0_0_0_a3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_data_0_LC_7_27_0 .C_ON=1'b0;
    defparam \my_uart.rx_data_0_LC_7_27_0 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_data_0_LC_7_27_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \my_uart.rx_data_0_LC_7_27_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1599),
            .lcout(LED_o_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2960),
            .ce(N__2063),
            .sr(_gnd_net_));
    defparam \my_uart.rx_data_7_LC_7_27_1 .C_ON=1'b0;
    defparam \my_uart.rx_data_7_LC_7_27_1 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_data_7_LC_7_27_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \my_uart.rx_data_7_LC_7_27_1  (
            .in0(N__3834),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(LED_o_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2960),
            .ce(N__2063),
            .sr(_gnd_net_));
    defparam \my_uart.rx_data_5_LC_7_27_2 .C_ON=1'b0;
    defparam \my_uart.rx_data_5_LC_7_27_2 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_data_5_LC_7_27_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \my_uart.rx_data_5_LC_7_27_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1662),
            .lcout(LED_o_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2960),
            .ce(N__2063),
            .sr(_gnd_net_));
    defparam \my_uart.rx_data_2_LC_7_27_3 .C_ON=1'b0;
    defparam \my_uart.rx_data_2_LC_7_27_3 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_data_2_LC_7_27_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \my_uart.rx_data_2_LC_7_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1641),
            .lcout(LED_o_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2960),
            .ce(N__2063),
            .sr(_gnd_net_));
    defparam \my_uart.rx_data_6_LC_7_27_4 .C_ON=1'b0;
    defparam \my_uart.rx_data_6_LC_7_27_4 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_data_6_LC_7_27_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \my_uart.rx_data_6_LC_7_27_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1683),
            .lcout(LED_o_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2960),
            .ce(N__2063),
            .sr(_gnd_net_));
    defparam \my_uart.rx_data_3_LC_7_27_5 .C_ON=1'b0;
    defparam \my_uart.rx_data_3_LC_7_27_5 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_data_3_LC_7_27_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \my_uart.rx_data_3_LC_7_27_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1560),
            .lcout(LED_o_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2960),
            .ce(N__2063),
            .sr(_gnd_net_));
    defparam \my_uart.rx_data_1_LC_7_27_6 .C_ON=1'b0;
    defparam \my_uart.rx_data_1_LC_7_27_6 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_data_1_LC_7_27_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \my_uart.rx_data_1_LC_7_27_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1620),
            .lcout(LED_o_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2960),
            .ce(N__2063),
            .sr(_gnd_net_));
    defparam \my_uart.rx_data_4_LC_7_27_7 .C_ON=1'b0;
    defparam \my_uart.rx_data_4_LC_7_27_7 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_data_4_LC_7_27_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \my_uart.rx_data_4_LC_7_27_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1578),
            .lcout(LED_o_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2960),
            .ce(N__2063),
            .sr(_gnd_net_));
    defparam \my_uart.rx_clk_divider_0_LC_9_25_0 .C_ON=1'b1;
    defparam \my_uart.rx_clk_divider_0_LC_9_25_0 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_clk_divider_0_LC_9_25_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \my_uart.rx_clk_divider_0_LC_9_25_0  (
            .in0(N__2681),
            .in1(N__1744),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\my_uart.rx_clk_dividerZ0Z_1 ),
            .ltout(),
            .carryin(bfn_9_25_0_),
            .carryout(\my_uart.rx_clk_divider_1_cry_0 ),
            .clk(N__2961),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_9_25_1 .C_ON=1'b1;
    defparam \my_uart.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_9_25_1 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_9_25_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \my_uart.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_9_25_1  (
            .in0(_gnd_net_),
            .in1(N__1711),
            .in2(N__2197),
            .in3(N__1549),
            .lcout(\my_uart.rx_clk_divider_1_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\my_uart.rx_clk_divider_1_cry_0 ),
            .carryout(\my_uart.rx_clk_divider_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_9_25_2 .C_ON=1'b1;
    defparam \my_uart.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_9_25_2 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_9_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \my_uart.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_9_25_2  (
            .in0(_gnd_net_),
            .in1(N__1900),
            .in2(N__2201),
            .in3(N__1546),
            .lcout(\my_uart.rx_clk_divider_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\my_uart.rx_clk_divider_1_cry_1 ),
            .carryout(\my_uart.rx_clk_divider_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_clk_divider_1_cry_2_THRU_LUT4_0_LC_9_25_3 .C_ON=1'b1;
    defparam \my_uart.rx_clk_divider_1_cry_2_THRU_LUT4_0_LC_9_25_3 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_clk_divider_1_cry_2_THRU_LUT4_0_LC_9_25_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \my_uart.rx_clk_divider_1_cry_2_THRU_LUT4_0_LC_9_25_3  (
            .in0(_gnd_net_),
            .in1(N__1783),
            .in2(N__2198),
            .in3(N__1543),
            .lcout(\my_uart.rx_clk_divider_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\my_uart.rx_clk_divider_1_cry_2 ),
            .carryout(\my_uart.rx_clk_divider_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_9_25_4 .C_ON=1'b1;
    defparam \my_uart.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_9_25_4 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_9_25_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \my_uart.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_9_25_4  (
            .in0(_gnd_net_),
            .in1(N__1827),
            .in2(N__2202),
            .in3(N__1765),
            .lcout(\my_uart.rx_clk_divider_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\my_uart.rx_clk_divider_1_cry_3 ),
            .carryout(\my_uart.rx_clk_divider_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_clk_divider_1_cry_4_THRU_LUT4_0_LC_9_25_5 .C_ON=1'b1;
    defparam \my_uart.rx_clk_divider_1_cry_4_THRU_LUT4_0_LC_9_25_5 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_clk_divider_1_cry_4_THRU_LUT4_0_LC_9_25_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \my_uart.rx_clk_divider_1_cry_4_THRU_LUT4_0_LC_9_25_5  (
            .in0(_gnd_net_),
            .in1(N__1849),
            .in2(N__2199),
            .in3(N__1762),
            .lcout(\my_uart.rx_clk_divider_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\my_uart.rx_clk_divider_1_cry_4 ),
            .carryout(\my_uart.rx_clk_divider_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_clk_divider_1_cry_5_THRU_LUT4_0_LC_9_25_6 .C_ON=1'b1;
    defparam \my_uart.rx_clk_divider_1_cry_5_THRU_LUT4_0_LC_9_25_6 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_clk_divider_1_cry_5_THRU_LUT4_0_LC_9_25_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \my_uart.rx_clk_divider_1_cry_5_THRU_LUT4_0_LC_9_25_6  (
            .in0(_gnd_net_),
            .in1(N__1804),
            .in2(N__2203),
            .in3(N__1759),
            .lcout(\my_uart.rx_clk_divider_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\my_uart.rx_clk_divider_1_cry_5 ),
            .carryout(\my_uart.rx_clk_divider_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_9_25_7 .C_ON=1'b1;
    defparam \my_uart.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_9_25_7 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_9_25_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \my_uart.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_9_25_7  (
            .in0(_gnd_net_),
            .in1(N__1933),
            .in2(N__2200),
            .in3(N__1756),
            .lcout(\my_uart.rx_clk_divider_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\my_uart.rx_clk_divider_1_cry_6 ),
            .carryout(\my_uart.rx_clk_divider_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_9_26_0 .C_ON=1'b1;
    defparam \my_uart.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_9_26_0 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_9_26_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \my_uart.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_9_26_0  (
            .in0(_gnd_net_),
            .in1(N__1962),
            .in2(N__2226),
            .in3(N__1753),
            .lcout(\my_uart.rx_clk_divider_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_9_26_0_),
            .carryout(\my_uart.rx_clk_divider_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_9_26_1 .C_ON=1'b1;
    defparam \my_uart.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_9_26_1 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_9_26_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \my_uart.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_9_26_1  (
            .in0(_gnd_net_),
            .in1(N__2220),
            .in2(N__2035),
            .in3(N__1750),
            .lcout(\my_uart.rx_clk_divider_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\my_uart.rx_clk_divider_1_cry_8 ),
            .carryout(\my_uart.rx_clk_divider_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_clk_divider_10_LC_9_26_2 .C_ON=1'b0;
    defparam \my_uart.rx_clk_divider_10_LC_9_26_2 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_clk_divider_10_LC_9_26_2 .LUT_INIT=16'b0010001000010001;
    LogicCell40 \my_uart.rx_clk_divider_10_LC_9_26_2  (
            .in0(N__1731),
            .in1(N__2688),
            .in2(_gnd_net_),
            .in3(N__1747),
            .lcout(\my_uart.rx_clk_dividerZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2963),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_clk_divider_RNIKT1U_10_LC_9_26_3 .C_ON=1'b0;
    defparam \my_uart.rx_clk_divider_RNIKT1U_10_LC_9_26_3 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_clk_divider_RNIKT1U_10_LC_9_26_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \my_uart.rx_clk_divider_RNIKT1U_10_LC_9_26_3  (
            .in0(N__1898),
            .in1(N__1743),
            .in2(N__1732),
            .in3(N__1709),
            .lcout(\my_uart.un1_rx_clk_divider_a_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_clk_divider_1_LC_9_26_4 .C_ON=1'b0;
    defparam \my_uart.rx_clk_divider_1_LC_9_26_4 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_clk_divider_1_LC_9_26_4 .LUT_INIT=16'b0000000010011001;
    LogicCell40 \my_uart.rx_clk_divider_1_LC_9_26_4  (
            .in0(N__1710),
            .in1(N__1717),
            .in2(_gnd_net_),
            .in3(N__2689),
            .lcout(\my_uart.rx_clk_dividerZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2963),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_clk_divider_8_LC_9_26_5 .C_ON=1'b0;
    defparam \my_uart.rx_clk_divider_8_LC_9_26_5 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_clk_divider_8_LC_9_26_5 .LUT_INIT=16'b1111111111111001;
    LogicCell40 \my_uart.rx_clk_divider_8_LC_9_26_5  (
            .in0(N__1963),
            .in1(N__1918),
            .in2(N__2701),
            .in3(N__2885),
            .lcout(\my_uart.rx_clk_dividerZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2963),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_clk_divider_9_LC_9_26_6 .C_ON=1'b0;
    defparam \my_uart.rx_clk_divider_9_LC_9_26_6 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_clk_divider_9_LC_9_26_6 .LUT_INIT=16'b0010001000010001;
    LogicCell40 \my_uart.rx_clk_divider_9_LC_9_26_6  (
            .in0(N__2033),
            .in1(N__2696),
            .in2(_gnd_net_),
            .in3(N__1912),
            .lcout(\my_uart.rx_clk_dividerZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2963),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_clk_divider_2_LC_9_26_7 .C_ON=1'b0;
    defparam \my_uart.rx_clk_divider_2_LC_9_26_7 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_clk_divider_2_LC_9_26_7 .LUT_INIT=16'b0000101000000101;
    LogicCell40 \my_uart.rx_clk_divider_2_LC_9_26_7  (
            .in0(N__1899),
            .in1(_gnd_net_),
            .in2(N__2700),
            .in3(N__1906),
            .lcout(\my_uart.rx_clk_dividerZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2963),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_clk_divider_3_LC_9_27_1 .C_ON=1'b0;
    defparam \my_uart.rx_clk_divider_3_LC_9_27_1 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_clk_divider_3_LC_9_27_1 .LUT_INIT=16'b1111111111111001;
    LogicCell40 \my_uart.rx_clk_divider_3_LC_9_27_1  (
            .in0(N__1779),
            .in1(N__1885),
            .in2(N__2699),
            .in3(N__2887),
            .lcout(\my_uart.rx_clk_dividerZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2965),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_clk_divider_4_LC_9_27_2 .C_ON=1'b0;
    defparam \my_uart.rx_clk_divider_4_LC_9_27_2 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_clk_divider_4_LC_9_27_2 .LUT_INIT=16'b1111111111101011;
    LogicCell40 \my_uart.rx_clk_divider_4_LC_9_27_2  (
            .in0(N__2888),
            .in1(N__1876),
            .in2(N__1828),
            .in3(N__2685),
            .lcout(\my_uart.rx_clk_dividerZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2965),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_clk_divider_6_LC_9_27_3 .C_ON=1'b0;
    defparam \my_uart.rx_clk_divider_6_LC_9_27_3 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_clk_divider_6_LC_9_27_3 .LUT_INIT=16'b0100010000010001;
    LogicCell40 \my_uart.rx_clk_divider_6_LC_9_27_3  (
            .in0(N__2687),
            .in1(N__1867),
            .in2(_gnd_net_),
            .in3(N__1799),
            .lcout(\my_uart.rx_clk_dividerZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2965),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_clk_divider_5_LC_9_27_4 .C_ON=1'b0;
    defparam \my_uart.rx_clk_divider_5_LC_9_27_4 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_clk_divider_5_LC_9_27_4 .LUT_INIT=16'b1111111011101111;
    LogicCell40 \my_uart.rx_clk_divider_5_LC_9_27_4  (
            .in0(N__2889),
            .in1(N__2686),
            .in2(N__1848),
            .in3(N__1858),
            .lcout(\my_uart.rx_clk_dividerZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2965),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_clk_divider_RNIIMPV_3_LC_9_27_6 .C_ON=1'b0;
    defparam \my_uart.rx_clk_divider_RNIIMPV_3_LC_9_27_6 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_clk_divider_RNIIMPV_3_LC_9_27_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \my_uart.rx_clk_divider_RNIIMPV_3_LC_9_27_6  (
            .in0(N__1841),
            .in1(N__1820),
            .in2(N__1803),
            .in3(N__1778),
            .lcout(\my_uart.un1_rx_clk_divider_a_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_10_24_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_10_24_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_10_24_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_10_24_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_RNO_5_2_LC_10_25_0 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_RNO_5_2_LC_10_25_0 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_RNO_5_2_LC_10_25_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \my_uart.rx_countdown_RNO_5_2_LC_10_25_0  (
            .in0(_gnd_net_),
            .in1(N__2419),
            .in2(_gnd_net_),
            .in3(N__2768),
            .lcout(\my_uart.rx_countdown_RNO_5Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_RNO_0_5_LC_10_25_1 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_RNO_0_5_LC_10_25_1 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_RNO_0_5_LC_10_25_1 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \my_uart.rx_countdown_RNO_0_5_LC_10_25_1  (
            .in0(N__3081),
            .in1(N__2537),
            .in2(N__2781),
            .in3(N__2864),
            .lcout(),
            .ltout(\my_uart.rx_countdown_8_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_5_LC_10_25_2 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_5_LC_10_25_2 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_countdown_5_LC_10_25_2 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \my_uart.rx_countdown_5_LC_10_25_2  (
            .in0(N__2677),
            .in1(_gnd_net_),
            .in2(N__1966),
            .in3(_gnd_net_),
            .lcout(\my_uart.rx_countdownZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2962),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_clk_divider_RNIF1TF_7_LC_10_25_3 .C_ON=1'b0;
    defparam \my_uart.rx_clk_divider_RNIF1TF_7_LC_10_25_3 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_clk_divider_RNIF1TF_7_LC_10_25_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \my_uart.rx_clk_divider_RNIF1TF_7_LC_10_25_3  (
            .in0(_gnd_net_),
            .in1(N__1961),
            .in2(_gnd_net_),
            .in3(N__1931),
            .lcout(\my_uart.un1_rx_clk_divider_a_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_RNO_6_2_LC_10_25_4 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_RNO_6_2_LC_10_25_4 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_RNO_6_2_LC_10_25_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \my_uart.rx_countdown_RNO_6_2_LC_10_25_4  (
            .in0(_gnd_net_),
            .in1(N__3080),
            .in2(_gnd_net_),
            .in3(N__3358),
            .lcout(),
            .ltout(\my_uart.rx_countdown_RNO_6Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_RNO_4_2_LC_10_25_5 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_RNO_4_2_LC_10_25_5 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_RNO_4_2_LC_10_25_5 .LUT_INIT=16'b0011111111011101;
    LogicCell40 \my_uart.rx_countdown_RNO_4_2_LC_10_25_5  (
            .in0(N__1948),
            .in1(N__2863),
            .in2(N__1942),
            .in3(N__3656),
            .lcout(\my_uart.rx_countdown_RNO_4Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_clk_divider_7_LC_10_25_6 .C_ON=1'b0;
    defparam \my_uart.rx_clk_divider_7_LC_10_25_6 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_clk_divider_7_LC_10_25_6 .LUT_INIT=16'b0000101000000101;
    LogicCell40 \my_uart.rx_clk_divider_7_LC_10_25_6  (
            .in0(N__1932),
            .in1(_gnd_net_),
            .in2(N__2698),
            .in3(N__1939),
            .lcout(\my_uart.rx_clk_dividerZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2962),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_RNIDTTP_2_LC_10_25_7 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_RNIDTTP_2_LC_10_25_7 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_RNIDTTP_2_LC_10_25_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \my_uart.rx_countdown_RNIDTTP_2_LC_10_25_7  (
            .in0(N__2318),
            .in1(N__2369),
            .in2(N__2496),
            .in3(N__3655),
            .lcout(\my_uart.g0_4_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_1_LC_10_26_1 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_1_LC_10_26_1 .SEQ_MODE=4'b1001;
    defparam \my_uart.rx_countdown_1_LC_10_26_1 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \my_uart.rx_countdown_1_LC_10_26_1  (
            .in0(N__2426),
            .in1(N__2552),
            .in2(N__2897),
            .in3(N__3361),
            .lcout(\my_uart.rx_countdownZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2964),
            .ce(),
            .sr(N__2697));
    defparam \my_uart.rx_countdown_RNO_0_2_LC_10_26_2 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_RNO_0_2_LC_10_26_2 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_RNO_0_2_LC_10_26_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \my_uart.rx_countdown_RNO_0_2_LC_10_26_2  (
            .in0(N__2367),
            .in1(N__2877),
            .in2(_gnd_net_),
            .in3(N__3188),
            .lcout(),
            .ltout(\my_uart.N_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_2_LC_10_26_3 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_2_LC_10_26_3 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_countdown_2_LC_10_26_3 .LUT_INIT=16'b1111111110101000;
    LogicCell40 \my_uart.rx_countdown_2_LC_10_26_3  (
            .in0(N__3727),
            .in1(N__2068),
            .in2(N__2044),
            .in3(N__2113),
            .lcout(\my_uart.rx_countdownZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2964),
            .ce(),
            .sr(N__2697));
    defparam \my_uart.rx_clk_divider_RNIU7NL2_9_LC_10_26_5 .C_ON=1'b0;
    defparam \my_uart.rx_clk_divider_RNIU7NL2_9_LC_10_26_5 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_clk_divider_RNIU7NL2_9_LC_10_26_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \my_uart.rx_clk_divider_RNIU7NL2_9_LC_10_26_5  (
            .in0(N__2041),
            .in1(N__2034),
            .in2(N__2011),
            .in3(N__2002),
            .lcout(\my_uart.un1_rx_clk_divider_a ),
            .ltout(\my_uart.un1_rx_clk_divider_a_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_RNIJ5KS3_5_LC_10_26_6 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_RNIJ5KS3_5_LC_10_26_6 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_RNIJ5KS3_5_LC_10_26_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \my_uart.rx_countdown_RNIJ5KS3_5_LC_10_26_6  (
            .in0(N__2776),
            .in1(N__1981),
            .in2(N__1993),
            .in3(N__2425),
            .lcout(\my_uart.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_RNIDTTP_0_2_LC_10_26_7 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_RNIDTTP_0_2_LC_10_26_7 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_RNIDTTP_0_2_LC_10_26_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \my_uart.rx_countdown_RNIDTTP_0_2_LC_10_26_7  (
            .in0(N__2305),
            .in1(N__2366),
            .in2(N__2488),
            .in3(N__3654),
            .lcout(\my_uart.g0_0_0_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNO_6_0_LC_10_27_0 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNO_6_0_LC_10_27_0 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNO_6_0_LC_10_27_0 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \my_uart.recv_state_RNO_6_0_LC_10_27_0  (
            .in0(N__3421),
            .in1(N__2242),
            .in2(N__3304),
            .in3(N__2778),
            .lcout(),
            .ltout(\my_uart.g0_6_a5_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNO_1_0_LC_10_27_1 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNO_1_0_LC_10_27_1 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNO_1_0_LC_10_27_1 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \my_uart.recv_state_RNO_1_0_LC_10_27_1  (
            .in0(N__2862),
            .in1(N__1972),
            .in2(N__1975),
            .in3(N__2092),
            .lcout(\my_uart.g0_6_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_4_LC_10_27_2 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_4_LC_10_27_2 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_countdown_4_LC_10_27_2 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \my_uart.rx_countdown_4_LC_10_27_2  (
            .in0(N__2131),
            .in1(_gnd_net_),
            .in2(N__2557),
            .in3(N__2633),
            .lcout(\my_uart.rx_countdownZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2966),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNO_5_0_LC_10_27_3 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNO_5_0_LC_10_27_3 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNO_5_0_LC_10_27_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \my_uart.recv_state_RNO_5_0_LC_10_27_3  (
            .in0(N__2368),
            .in1(N__2312),
            .in2(N__2489),
            .in3(N__2420),
            .lcout(\my_uart.g0_6_a5_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_3_LC_10_27_4 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_3_LC_10_27_4 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_countdown_3_LC_10_27_4 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \my_uart.rx_countdown_3_LC_10_27_4  (
            .in0(N__2553),
            .in1(N__2632),
            .in2(_gnd_net_),
            .in3(N__2107),
            .lcout(\my_uart.rx_countdownZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2966),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_RNINCD63_4_LC_10_27_5 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_RNINCD63_4_LC_10_27_5 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_RNINCD63_4_LC_10_27_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \my_uart.rx_countdown_RNINCD63_4_LC_10_27_5  (
            .in0(N__2480),
            .in1(_gnd_net_),
            .in2(N__2890),
            .in3(N__3130),
            .lcout(\my_uart.rx_countdown_3_4 ),
            .ltout(\my_uart.rx_countdown_3_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_RNO_2_2_LC_10_27_6 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_RNO_2_2_LC_10_27_6 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_RNO_2_2_LC_10_27_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \my_uart.rx_countdown_RNO_2_2_LC_10_27_6  (
            .in0(N__2098),
            .in1(N__2106),
            .in2(N__2125),
            .in3(N__2122),
            .lcout(\my_uart.N_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_RNIK53C3_3_LC_10_27_7 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_RNIK53C3_3_LC_10_27_7 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_RNIK53C3_3_LC_10_27_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \my_uart.rx_countdown_RNIK53C3_3_LC_10_27_7  (
            .in0(N__2858),
            .in1(N__2313),
            .in2(_gnd_net_),
            .in3(N__3714),
            .lcout(\my_uart.rx_countdown_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_RNO_3_2_LC_10_28_2 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_RNO_3_2_LC_10_28_2 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_RNO_3_2_LC_10_28_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \my_uart.rx_countdown_RNO_3_2_LC_10_28_2  (
            .in0(N__3245),
            .in1(N__3420),
            .in2(N__3832),
            .in3(N__3560),
            .lcout(\my_uart.G_14_0_a3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNO_4_0_LC_10_28_6 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNO_4_0_LC_10_28_6 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNO_4_0_LC_10_28_6 .LUT_INIT=16'b0111011100000001;
    LogicCell40 \my_uart.recv_state_RNO_4_0_LC_10_28_6  (
            .in0(N__3244),
            .in1(N__3419),
            .in2(N__3831),
            .in3(N__3559),
            .lcout(\my_uart.g0_6_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_RNIEMHI6_2_LC_11_25_0 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_RNIEMHI6_2_LC_11_25_0 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_RNIEMHI6_2_LC_11_25_0 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \my_uart.rx_countdown_RNIEMHI6_2_LC_11_25_0  (
            .in0(N__2871),
            .in1(N__2248),
            .in2(N__2086),
            .in3(N__2260),
            .lcout(),
            .ltout(\my_uart.rx_countdown20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNIG81F7_1_LC_11_25_1 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNIG81F7_1_LC_11_25_1 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNIG81F7_1_LC_11_25_1 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \my_uart.recv_state_RNIG81F7_1_LC_11_25_1  (
            .in0(N__2074),
            .in1(_gnd_net_),
            .in2(N__2077),
            .in3(N__2254),
            .lcout(\my_uart.un1_rx_data_0_sqmuxa_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNIOPND_1_1_LC_11_25_2 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNIOPND_1_1_LC_11_25_2 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNIOPND_1_1_LC_11_25_2 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \my_uart.recv_state_RNIOPND_1_1_LC_11_25_2  (
            .in0(N__3540),
            .in1(_gnd_net_),
            .in2(N__3459),
            .in3(N__3299),
            .lcout(\my_uart.un1_recv_state_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNIOPND_1_LC_11_25_3 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNIOPND_1_LC_11_25_3 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNIOPND_1_LC_11_25_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \my_uart.recv_state_RNIOPND_1_LC_11_25_3  (
            .in0(N__3297),
            .in1(N__3447),
            .in2(_gnd_net_),
            .in3(N__3538),
            .lcout(\my_uart.un1_recv_state_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_RNIH36N1_0_0_LC_11_25_4 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_RNIH36N1_0_0_LC_11_25_4 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_RNIH36N1_0_0_LC_11_25_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \my_uart.rx_countdown_RNIH36N1_0_0_LC_11_25_4  (
            .in0(N__3189),
            .in1(N__3647),
            .in2(N__3362),
            .in3(N__3710),
            .lcout(),
            .ltout(\my_uart.g0_4_a3_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_RNIRGTL2_0_LC_11_25_5 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_RNIRGTL2_0_LC_11_25_5 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_RNIRGTL2_0_LC_11_25_5 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \my_uart.rx_countdown_RNIRGTL2_0_LC_11_25_5  (
            .in0(_gnd_net_),
            .in1(N__3124),
            .in2(N__2263),
            .in3(N__3082),
            .lcout(\my_uart.g0_4_a3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNIAONE_1_LC_11_25_6 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNIAONE_1_LC_11_25_6 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNIAONE_1_LC_11_25_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \my_uart.recv_state_RNIAONE_1_LC_11_25_6  (
            .in0(N__3539),
            .in1(N__3806),
            .in2(N__3458),
            .in3(N__3298),
            .lcout(\my_uart.recv_state_0_sqmuxa_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_RNI80VC_5_LC_11_25_7 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_RNI80VC_5_LC_11_25_7 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_RNI80VC_5_LC_11_25_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \my_uart.rx_countdown_RNI80VC_5_LC_11_25_7  (
            .in0(_gnd_net_),
            .in1(N__2772),
            .in2(_gnd_net_),
            .in3(N__2421),
            .lcout(\my_uart.g0_4_a3_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNO_8_0_LC_11_26_0 .C_ON=1'b1;
    defparam \my_uart.recv_state_RNO_8_0_LC_11_26_0 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNO_8_0_LC_11_26_0 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \my_uart.recv_state_RNO_8_0_LC_11_26_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3662),
            .in3(N__3516),
            .lcout(\my_uart.g0_6_a5_1_0 ),
            .ltout(),
            .carryin(bfn_11_26_0_),
            .carryout(\my_uart.rx_countdown_3_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_3_cry_0_s1_c_RNIE18B_LC_11_26_1 .C_ON=1'b1;
    defparam \my_uart.rx_countdown_3_cry_0_s1_c_RNIE18B_LC_11_26_1 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_3_cry_0_s1_c_RNIE18B_LC_11_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \my_uart.rx_countdown_3_cry_0_s1_c_RNIE18B_LC_11_26_1  (
            .in0(_gnd_net_),
            .in1(N__2209),
            .in2(N__2427),
            .in3(N__2236),
            .lcout(\my_uart.rx_countdown_3_s1_1 ),
            .ltout(),
            .carryin(\my_uart.rx_countdown_3_cry_0_s1 ),
            .carryout(\my_uart.rx_countdown_3_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_3_cry_1_s1_c_RNIG7IL_LC_11_26_2 .C_ON=1'b1;
    defparam \my_uart.rx_countdown_3_cry_1_s1_c_RNIG7IL_LC_11_26_2 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_3_cry_1_s1_c_RNIG7IL_LC_11_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \my_uart.rx_countdown_3_cry_1_s1_c_RNIG7IL_LC_11_26_2  (
            .in0(_gnd_net_),
            .in1(N__2221),
            .in2(N__2370),
            .in3(N__2233),
            .lcout(\my_uart.rx_countdown_3_s1_2 ),
            .ltout(),
            .carryin(\my_uart.rx_countdown_3_cry_1_s1 ),
            .carryout(\my_uart.rx_countdown_3_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_3_cry_2_s1_c_RNIIDSF_LC_11_26_3 .C_ON=1'b1;
    defparam \my_uart.rx_countdown_3_cry_2_s1_c_RNIIDSF_LC_11_26_3 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_3_cry_2_s1_c_RNIIDSF_LC_11_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \my_uart.rx_countdown_3_cry_2_s1_c_RNIIDSF_LC_11_26_3  (
            .in0(_gnd_net_),
            .in1(N__2304),
            .in2(N__2227),
            .in3(N__2230),
            .lcout(\my_uart.rx_countdown_3_s1_3 ),
            .ltout(),
            .carryin(\my_uart.rx_countdown_3_cry_2_s1 ),
            .carryout(\my_uart.rx_countdown_3_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_3_cry_3_s1_c_RNIKJ6A_LC_11_26_4 .C_ON=1'b1;
    defparam \my_uart.rx_countdown_3_cry_3_s1_c_RNIKJ6A_LC_11_26_4 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_3_cry_3_s1_c_RNIKJ6A_LC_11_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \my_uart.rx_countdown_3_cry_3_s1_c_RNIKJ6A_LC_11_26_4  (
            .in0(_gnd_net_),
            .in1(N__2225),
            .in2(N__2484),
            .in3(N__2563),
            .lcout(\my_uart.rx_countdown_3_s1_4 ),
            .ltout(),
            .carryin(\my_uart.rx_countdown_3_cry_3_s1 ),
            .carryout(\my_uart.rx_countdown_3_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_3_cry_4_s1_c_RNIMPGK_LC_11_26_5 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_3_cry_4_s1_c_RNIMPGK_LC_11_26_5 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_3_cry_4_s1_c_RNIMPGK_LC_11_26_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \my_uart.rx_countdown_3_cry_4_s1_c_RNIMPGK_LC_11_26_5  (
            .in0(_gnd_net_),
            .in1(N__2777),
            .in2(_gnd_net_),
            .in3(N__2560),
            .lcout(\my_uart.rx_countdown_3_s1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_0_LC_11_26_6 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_0_LC_11_26_6 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_countdown_0_LC_11_26_6 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \my_uart.rx_countdown_0_LC_11_26_6  (
            .in0(N__3646),
            .in1(N__2538),
            .in2(N__2676),
            .in3(N__2886),
            .lcout(\my_uart.rx_countdownZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2967),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_bits_remaining_RNO_6_3_LC_11_26_7 .C_ON=1'b0;
    defparam \my_uart.rx_bits_remaining_RNO_6_3_LC_11_26_7 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_bits_remaining_RNO_6_3_LC_11_26_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \my_uart.rx_bits_remaining_RNO_6_3_LC_11_26_7  (
            .in0(N__3178),
            .in1(N__3645),
            .in2(N__3363),
            .in3(N__3709),
            .lcout(\my_uart.g0_0_0_a3_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNO_0_1_LC_11_27_0 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNO_0_1_LC_11_27_0 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNO_0_1_LC_11_27_0 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \my_uart.recv_state_RNO_0_1_LC_11_27_0  (
            .in0(N__3586),
            .in1(N__2881),
            .in2(N__2506),
            .in3(N__2716),
            .lcout(),
            .ltout(\my_uart.N_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_1_LC_11_27_1 .C_ON=1'b0;
    defparam \my_uart.recv_state_1_LC_11_27_1 .SEQ_MODE=4'b1000;
    defparam \my_uart.recv_state_1_LC_11_27_1 .LUT_INIT=16'b0001110111000000;
    LogicCell40 \my_uart.recv_state_1_LC_11_27_1  (
            .in0(N__3530),
            .in1(N__3282),
            .in2(N__2509),
            .in3(N__3440),
            .lcout(N_18_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2969),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNO_4_1_LC_11_27_2 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNO_4_1_LC_11_27_2 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNO_4_1_LC_11_27_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \my_uart.recv_state_RNO_4_1_LC_11_27_2  (
            .in0(N__2470),
            .in1(N__2314),
            .in2(_gnd_net_),
            .in3(N__2361),
            .lcout(\my_uart.N_22_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNO_1_1_LC_11_27_3 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNO_1_1_LC_11_27_3 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNO_1_1_LC_11_27_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \my_uart.recv_state_RNO_1_1_LC_11_27_3  (
            .in0(N__2418),
            .in1(N__2779),
            .in2(N__3556),
            .in3(N__3659),
            .lcout(\my_uart.N_18_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNO_4_2_LC_11_27_4 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNO_4_2_LC_11_27_4 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNO_4_2_LC_11_27_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \my_uart.recv_state_RNO_4_2_LC_11_27_4  (
            .in0(N__2469),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2417),
            .lcout(),
            .ltout(\my_uart.m10_e_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNO_2_2_LC_11_27_5 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNO_2_2_LC_11_27_5 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNO_2_2_LC_11_27_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \my_uart.recv_state_RNO_2_2_LC_11_27_5  (
            .in0(N__2362),
            .in1(N__2322),
            .in2(N__2266),
            .in3(N__2780),
            .lcout(\my_uart.m10_e_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNO_5_1_LC_11_27_6 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNO_5_1_LC_11_27_6 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNO_5_1_LC_11_27_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \my_uart.recv_state_RNO_5_1_LC_11_27_6  (
            .in0(N__3122),
            .in1(N__3186),
            .in2(_gnd_net_),
            .in3(N__3715),
            .lcout(),
            .ltout(\my_uart.N_23_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNO_3_1_LC_11_27_7 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNO_3_1_LC_11_27_7 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNO_3_1_LC_11_27_7 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \my_uart.recv_state_RNO_3_1_LC_11_27_7  (
            .in0(N__3833),
            .in1(N__2725),
            .in2(N__2719),
            .in3(N__3660),
            .lcout(\my_uart.m7_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNO_0_0_LC_11_28_0 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNO_0_0_LC_11_28_0 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNO_0_0_LC_11_28_0 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \my_uart.recv_state_RNO_0_0_LC_11_28_0  (
            .in0(N__2710),
            .in1(N__2898),
            .in2(N__3142),
            .in3(N__3673),
            .lcout(),
            .ltout(\my_uart.un1_rx_clk_divider28_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_0_LC_11_28_1 .C_ON=1'b0;
    defparam \my_uart.recv_state_0_LC_11_28_1 .SEQ_MODE=4'b1000;
    defparam \my_uart.recv_state_0_LC_11_28_1 .LUT_INIT=16'b1111101000111010;
    LogicCell40 \my_uart.recv_state_0_LC_11_28_1  (
            .in0(N__3274),
            .in1(N__2599),
            .in2(N__2704),
            .in3(N__3466),
            .lcout(my_uart_recv_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2971),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNIAONE_0_1_LC_11_28_3 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNIAONE_0_1_LC_11_28_3 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNIAONE_0_1_LC_11_28_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \my_uart.recv_state_RNIAONE_0_1_LC_11_28_3  (
            .in0(N__3272),
            .in1(N__3437),
            .in2(N__3829),
            .in3(N__3554),
            .lcout(\my_uart.rx_clk_divider_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_cnst_2_0__m6_0_18_0_LC_11_28_5 .C_ON=1'b0;
    defparam \my_uart.recv_state_cnst_2_0__m6_0_18_0_LC_11_28_5 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_cnst_2_0__m6_0_18_0_LC_11_28_5 .LUT_INIT=16'b1111011111000110;
    LogicCell40 \my_uart.recv_state_cnst_2_0__m6_0_18_0_LC_11_28_5  (
            .in0(N__3273),
            .in1(N__3438),
            .in2(N__3830),
            .in3(N__3555),
            .lcout(\my_uart.m6_0_18_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_cnst_2_0__m6_0_18_a4_1_2_LC_12_25_0 .C_ON=1'b0;
    defparam \my_uart.recv_state_cnst_2_0__m6_0_18_a4_1_2_LC_12_25_0 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_cnst_2_0__m6_0_18_a4_1_2_LC_12_25_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \my_uart.recv_state_cnst_2_0__m6_0_18_a4_1_2_LC_12_25_0  (
            .in0(N__2993),
            .in1(N__3035),
            .in2(N__2593),
            .in3(N__3022),
            .lcout(\my_uart.m6_0_18_a4_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_bits_remaining_1_LC_12_25_1 .C_ON=1'b0;
    defparam \my_uart.rx_bits_remaining_1_LC_12_25_1 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_bits_remaining_1_LC_12_25_1 .LUT_INIT=16'b0000000010100101;
    LogicCell40 \my_uart.rx_bits_remaining_1_LC_12_25_1  (
            .in0(N__3025),
            .in1(_gnd_net_),
            .in2(N__3040),
            .in3(N__3302),
            .lcout(\my_uart.rx_bits_remainingZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2968),
            .ce(N__2980),
            .sr(_gnd_net_));
    defparam \my_uart.rx_bits_remaining_0_LC_12_25_3 .C_ON=1'b0;
    defparam \my_uart.rx_bits_remaining_0_LC_12_25_3 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_bits_remaining_0_LC_12_25_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \my_uart.rx_bits_remaining_0_LC_12_25_3  (
            .in0(N__3024),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3301),
            .lcout(\my_uart.rx_bits_remainingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2968),
            .ce(N__2980),
            .sr(_gnd_net_));
    defparam \my_uart.rx_bits_remaining_RNINFUH_1_LC_12_25_4 .C_ON=1'b0;
    defparam \my_uart.rx_bits_remaining_RNINFUH_1_LC_12_25_4 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_bits_remaining_RNINFUH_1_LC_12_25_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \my_uart.rx_bits_remaining_RNINFUH_1_LC_12_25_4  (
            .in0(_gnd_net_),
            .in1(N__3036),
            .in2(_gnd_net_),
            .in3(N__3023),
            .lcout(\my_uart.CO1_i ),
            .ltout(\my_uart.CO1_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_bits_remaining_2_LC_12_25_5 .C_ON=1'b0;
    defparam \my_uart.rx_bits_remaining_2_LC_12_25_5 .SEQ_MODE=4'b1000;
    defparam \my_uart.rx_bits_remaining_2_LC_12_25_5 .LUT_INIT=16'b0000000000111100;
    LogicCell40 \my_uart.rx_bits_remaining_2_LC_12_25_5  (
            .in0(_gnd_net_),
            .in1(N__2994),
            .in2(N__3001),
            .in3(N__3303),
            .lcout(\my_uart.rx_bits_remainingZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2968),
            .ce(N__2980),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_2_LC_12_26_0 .C_ON=1'b0;
    defparam \my_uart.recv_state_2_LC_12_26_0 .SEQ_MODE=4'b1000;
    defparam \my_uart.recv_state_2_LC_12_26_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \my_uart.recv_state_2_LC_12_26_0  (
            .in0(N__2788),
            .in1(N__2920),
            .in2(_gnd_net_),
            .in3(N__3661),
            .lcout(my_uart_recv_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2970),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNO_5_2_LC_12_26_1 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNO_5_2_LC_12_26_1 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNO_5_2_LC_12_26_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \my_uart.recv_state_RNO_5_2_LC_12_26_1  (
            .in0(_gnd_net_),
            .in1(N__3354),
            .in2(_gnd_net_),
            .in3(N__3185),
            .lcout(),
            .ltout(\my_uart.m15_e_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNO_3_2_LC_12_26_2 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNO_3_2_LC_12_26_2 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNO_3_2_LC_12_26_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \my_uart.recv_state_RNO_3_2_LC_12_26_2  (
            .in0(N__3131),
            .in1(N__3089),
            .in2(N__2926),
            .in3(N__3716),
            .lcout(),
            .ltout(\my_uart.m15_e_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNO_1_2_LC_12_26_3 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNO_1_2_LC_12_26_3 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNO_1_2_LC_12_26_3 .LUT_INIT=16'b0101110011001100;
    LogicCell40 \my_uart.recv_state_RNO_1_2_LC_12_26_3  (
            .in0(N__3736),
            .in1(N__2914),
            .in2(N__2923),
            .in3(N__2896),
            .lcout(\my_uart.N_28_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNIOPND_0_1_LC_12_26_4 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNIOPND_0_1_LC_12_26_4 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNIOPND_0_1_LC_12_26_4 .LUT_INIT=16'b0100010011111111;
    LogicCell40 \my_uart.recv_state_RNIOPND_0_1_LC_12_26_4  (
            .in0(N__3286),
            .in1(N__3423),
            .in2(_gnd_net_),
            .in3(N__3531),
            .lcout(\my_uart.N_19_mux_0 ),
            .ltout(\my_uart.N_19_mux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNO_0_2_LC_12_26_5 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNO_0_2_LC_12_26_5 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNO_0_2_LC_12_26_5 .LUT_INIT=16'b1111000001110100;
    LogicCell40 \my_uart.recv_state_RNO_0_2_LC_12_26_5  (
            .in0(N__3735),
            .in1(N__2908),
            .in2(N__2902),
            .in3(N__2895),
            .lcout(\my_uart.N_27_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RS232_RX_i_ibuf_RNIAONE_LC_12_26_6.C_ON=1'b0;
    defparam RS232_RX_i_ibuf_RNIAONE_LC_12_26_6.SEQ_MODE=4'b0000;
    defparam RS232_RX_i_ibuf_RNIAONE_LC_12_26_6.LUT_INIT=16'b1010101010101000;
    LogicCell40 RS232_RX_i_ibuf_RNIAONE_LC_12_26_6 (
            .in0(N__3287),
            .in1(N__3422),
            .in2(N__3828),
            .in3(N__3532),
            .lcout(N_20_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.rx_countdown_RNO_1_2_LC_12_26_7 .C_ON=1'b0;
    defparam \my_uart.rx_countdown_RNO_1_2_LC_12_26_7 .SEQ_MODE=4'b0000;
    defparam \my_uart.rx_countdown_RNO_1_2_LC_12_26_7 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \my_uart.rx_countdown_RNO_1_2_LC_12_26_7  (
            .in0(N__3533),
            .in1(N__3288),
            .in2(_gnd_net_),
            .in3(N__3439),
            .lcout(\my_uart.N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNO_3_0_LC_12_27_0 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNO_3_0_LC_12_27_0 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNO_3_0_LC_12_27_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \my_uart.recv_state_RNO_3_0_LC_12_27_0  (
            .in0(N__3658),
            .in1(N__3046),
            .in2(N__3558),
            .in3(N__3717),
            .lcout(\my_uart.g0_6_a5_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNO_2_1_LC_12_27_3 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNO_2_1_LC_12_27_3 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNO_2_1_LC_12_27_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \my_uart.recv_state_RNO_2_1_LC_12_27_3  (
            .in0(N__3088),
            .in1(N__3359),
            .in2(N__3557),
            .in3(N__3657),
            .lcout(\my_uart.N_19_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_cnst_2_0__m6_0_18_a4_1_LC_12_27_4 .C_ON=1'b0;
    defparam \my_uart.recv_state_cnst_2_0__m6_0_18_a4_1_LC_12_27_4 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_cnst_2_0__m6_0_18_a4_1_LC_12_27_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \my_uart.recv_state_cnst_2_0__m6_0_18_a4_1_LC_12_27_4  (
            .in0(N__3580),
            .in1(N__3271),
            .in2(_gnd_net_),
            .in3(N__3537),
            .lcout(\my_uart.N_217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNO_2_0_LC_12_27_5 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNO_2_0_LC_12_27_5 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNO_2_0_LC_12_27_5 .LUT_INIT=16'b0000000000110010;
    LogicCell40 \my_uart.recv_state_RNO_2_0_LC_12_27_5  (
            .in0(N__3436),
            .in1(N__3360),
            .in2(N__3300),
            .in3(N__3187),
            .lcout(\my_uart.g0_6_a5_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \my_uart.recv_state_RNO_7_0_LC_12_27_7 .C_ON=1'b0;
    defparam \my_uart.recv_state_RNO_7_0_LC_12_27_7 .SEQ_MODE=4'b0000;
    defparam \my_uart.recv_state_RNO_7_0_LC_12_27_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \my_uart.recv_state_RNO_7_0_LC_12_27_7  (
            .in0(_gnd_net_),
            .in1(N__3123),
            .in2(_gnd_net_),
            .in3(N__3079),
            .lcout(\my_uart.g0_6_a5_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // uart_top
